��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����`��B�㓪F:��ew���@�C�k�.U6�vά1�xrl9��Sr?$R�t��M��~3pwd��<�i��w_�)4ޟo$#)����4F�1s[�p;��Q�!����7�5G��Ξ@��/6����Q�&�$G��Fs���K�+������;V�P���l��X�g�rNR�;hVC��D}�LX���J�lq@Á]��d��择+I@��g�&�Nj�{q��"H_X�&Gbr��	��Q���=c�dG�	Wyp$MR�DP;`��|N�έ�����#m-�L�eBB��;�P���aY��	X;Pvi�+���L���5�f���k��"ƈ��^���(�a�R[��J��ksD�0�,;S<-t���{r�kg��f����A���7�H)7��@l�y�s_�'�5�+!�G>vo9���&��)�5u��jE���	���6-,;0g��݉��%r��1L�����X��H��X������~�d����/� ���k��k(7⅚z^�y���-��b�KiQ�,I�WDƎ�,�PS<-�tE[��f����	ԘR%E�0T�s-��{2Ł�z[nt����)�&�:�ζ<��+4�%��L��S��w��h�z� ��'�>�|�z���t����;�dT�T�&JM�B��� ���۞Pb.�A�!A��_sǯ1Z,��e�QI�$��Úly�햾�E��4e�O��sTp-.#sq�I�y�s���ww��̰����!Ƙ�0
�܆4 ��P �qC1$�J��R)�$��Q�����3u�8��BZ�J%�?Lu�\���d$	6��&��p�=� u�e͟\K�����֐�pV�#]�R�c�.���;���4���T���W�U��2k��Шo��[L���0�ӳ�����(���Q"˽������,/M��D)�щ��^�KO{���.Э4Z�y]�V-��!�� �7�'
��/�k֖�0�F%����x��l% J�8��>*��N)_�\µ�d'�#E~��7��|8��l�'�`upգj���PVm/�5Hl*����JFN�q=��A���wV}���"��o�@�S�D�J��F�K����>�H�  ��6�ކ���"� �|�$��ݚf��[�~ �Ge)��"�/�K�+�|��W�l9�r�2��[�P�eg����\�yn��<��\��=��Åˉ��Ö;�w�ϬWO�]�G��&ô*�!)�ޕ��`�&]�J/6�����f
�9[~�9/&W���B�q�p5��.e�cq�F����2uP��p�\��&7��1�ڄ�J5)�伶^��vQ�\rU����w6���>�*�ɯ�^כ��M��z���b��H�E�V3 �Cf&��j���+86_D���Q��k���1��(2�j�Z"k6�i�N�|�T���[1V �K�هVs�-v�1�:��ᙢ���m��U2�K���)yr�W�����@F~�yw��	���G4�`]R��>wAgf�o��[���]Y����xt���9�I:�д���5�Ø�����rCZ��>K	���<D�C��c�B6�u�f�T砝�[�*avr����af2A~j�:���ڎѻP�Xl�zɁ��"BL�;�5�ͩ;��7�V���UP]��-9�h�$1����3�{@o�cL/�^��p�^���E<�>$�l\�t���&H�^�^t'{_����jN')t����0>j���RM'h�����|P����aY�\�,��O9ܶM��_��M_���W���&B\�#���{Z��8d/H�W�s͇�'�� ��tl=�De-�L�׆t��k�8��(���Ą�����C�H_ӇG2�C*я�`����|F��9K=Yv�T��MﻓP3qۃ��#��i�r-�^��Cw�oؾ��Z�>��� a�����ǯ�i�qm/"����ݿ��Ǐ�����4(�+��a�_H�'�KB/�e��*]N�T�ɡ�2�܁�jS��؂����^o�I
?f���)ȉ{���+��<e��$Y�]⽾@�W��)O�r�\���!��sF;Ow��b��5.0.���`�#w��E�t�)��Q��Jx~,!9�T�� ������6]P<���i����	R=$�x�N�j�ǎy������┐_�.�Si�3��(��B���2�� s����R��x�&�2����^y5iNq:=�'�J��d���(�TT�.�u �2����1<g��c�#%�X��5�[]L	!��w�IjF�z���z�g&��w��()�l�$����3S@���%] �<���5�c�Q[O�m�#n2�����k|Q���8:)�n��T�6�}��
�-�dN�`<��t��SC�Ο���^�/t��;�j)�4n˜�s������_���Ð,���ꤙc�F�%�|�����<<s:{H�C��۷[�f<��A��[u����ਛ>d���R�{j]��+s�����Ck�[���{��o�"��w}�q-�r0\x@`�M�+�R�BAW^�:Ԟ�S��s�=���/f-u��|
=FIL8K^��b�TB�����无bU����On�DB��q<@�jv�wd ~t�ΟF���IX���k���_�i�ᆄ��i�����g�!3�+1QyM���G�-��#�F���QAAM�Q4����/�T�� ��r��K� ��^%ב̪�y���F����W�V���YrƉv�J{0�C�|�K�\��ue�'��fzU��2*�.�ay$-q�?�r��U0��A%�3�ԟ�}&�r )���������k^)�T�T��x�%��s}{7�>���(݃p�򯘅�I�S�Bo�[\a����H�����3L+��~%�Ͱ��\u�a� �ށ�b����pY^��uv#��������eM���®�UMP���ܽ�1��/��s���_��t���JY9��B7)�YS�`4.,<��prl��+�f��(�E-X��C�~���k�aY�gN�H��R� /�㶒@��с)�� 	���+IcC���im����,��FS��`�A���ܗ�P���ƿ���*�����������V�#���w&Wig~���[�$�� ��|:r���)�
�ל֪"PC��J� ˇl3�*���i�� y��;S$l�������c�6bV5��! W�+&��+d�9��(�e�UM�
;D����%���\��I`�6u_�NG��ˈ�ip�4��W�D����S��sk��'���9$N-��W��>Ѣ	��z�/�����q�sBJ������]U�%��G�|kn�4�lLN��dY0�Yh�Y߅iK��nMpD�fP\��YS�Jׂ���])�T�c�����P�`�f���iƹ��4-�q��h��#J���
�"�h��<U��׏���9t��f�E�=�=��l���&ސ���IU�]Rb�^�ᖈ<AWBO:��z"57X�cNa�K�V�I�	�9I�'�":���lrW̎rP��_)��x�U�`�F�y'��J�+�kRCNN����i�R1�X́$�6��T��aL΢����0�:sy�e����Ϻ)a8�6�kf������E�m��Lg"f���TW�S�c�#g&��x���c,�o���G��H�؟����*i�'k�[I)����x&V4:J��2ຩ��0̓����j%9l���!��3ZN�B�i%�$jA~&���q�<s��mB�ׇ)���F�k�u �eO~�0��62x��T���7��`2�u�Ƞ����x%�яPX�˒<�����>�L�-bl J*��w�F?�6�0\%/����]n�Eda�[Q��c3q7@�ɸ�q`�|r�Hr����4���Q�HH{�>�{�������(M���r���#S��l�i����7�گ�\��W�7��Yd�z$� h�[d�D��[4�'�ʼӪA�S>L ����h�_�uj*8\8y� Q��{}��v�t����C��e�X��("�;��Mc��1�#�~Z�*�VKJ|���t��NU+6&�:9�-&+
��}�PmvmH��ʤ����V�Qvp_6�\�7���O��f���Z�q�!&4e�1�v��ZL�NI�b���`�?ڣ�(�` ���K�_�?G~���'�8�r���8����ޏ�	� ��C]�tsU��D�3h��7}+9��~��W/��X�BI�y����J��4wdMG�,I7A���<X;�}�=���|�5�W��U�s��R����:��_K��%t����{�o�+�1h�x��7/g���]�I@ۈw�p����u�s��c��g�  j_��ޔ �U�6*���_n
z�H�}T`�(�:K�-�2 ��\B���e�y����-����:����U5I�s'};���?#+X�3u9�	@r�s��Z.�qor�a�K\���|!�ic���y�|1�z���v�-��$D�9�QT�?^�]��cg91��X����$ܤewb�k�{�f�E�ߩ�3�A��p̝3u���g�*u\��5��E)�ìZU���Lo��)�<���\�������x���?<b��Zm�?�v������W桊�qˎ7�1ח���͆���h_���${CBH�f�+�үƊ�h�� ��M��ܺ�y�z���*���i	ž�u�(�D&p����i��:!���ZÁQ�����;{�ҕsN&��D�4X�M�P]�n���r ���32��4K@�%E%����}��)3�$%³��ItLji�F�F��ٗ��� ���Y;����ȧ'k����bX+,���=c?��9����&�Fֵ͍}�{=:�?/��F�).��C��:���{�5�Eut�S��.��_m73��|�u��.3��E�7Q�l���%뮟�
�"����Ǘ�M��k����w�[Fm���͑�<�/���B���\�h}���dV�t�14d�<���@b�R���vT�
x%;IN��z��f�������m*ZOs�{U���h}����f`��v�Ev���ǖ,*Eap���π��C�ǜt�h�p��>�7�G�`mA���x�bt���}�g���S����h�v�^�zC|Ҳ ����������@�h���3[�� �ȋJ�1��u4���LTLVq*�d�ŽaB�d��'~���FS�����w>OK�I}�#�](�~�E˶��VgJAar�k�0��0�� ��]a3����Ķ8	X(�,�%�gX|k�E�i�������7
J��!`�"8����lf#�l>��0���;X����_f25xG).���z� :�!���}
қ�3*�Ȱ@m�Dh�M���U�-qJl�&h��a�����m%3�~uw9��N�̑S~�4�خY�!Psd$�U�L>�j��Y��Xjgw�ja�C�/ޓլUjpT�	��ǘP�a�,�<D ��.<��O�gGy'�)���<��N!��־L�*r�X˰���uss�I�t�=����hGho�
���T�^`���@�h�}kz�VRs+}{��Zݝ-����LZ`��Tq��������)ޟјz��C/� ��������-�tAJW��JP��~�>}�����+���"7D���N���b]���+(R
n��c@sQ�����X%�1�-媷/��Fb+�"1
w�`�p��'h���1��)�;��fq4b�d�[|�����_�J*:��������k�9��nfI/,����vm7π��M��ǭ�#���V"���E��x�҉������P���J��E^S�2���Sn�Eg���À_Xs���i7����l�E&��,�fu����m��p躹�����f�;���5@�Pi"AE���F*B�C}Bs]2�\��gH�S���5e�B/u�߃��J�Ucy�^H9�?�/ �@���+��_zZ_@�����ψ��87'Y�֙�ZM�W��Bd�?�Ǖ��D�u������J1(Z���V�qo.R�z�[:�y�R;z6/�A�w��p�P��|.�]�x�0�����w���]�e���.K5�ǂ�(�G��?.E�[g�����_Iv5 a��L`�8͢���s!�@`���r����T�3dn��󠪞�mhǕ9Kս�Nw?�y�������{pQ�c@��ù]-N�K⊬�|n��h)>[���-<	���;;���ގ��K�
���|=�{v��+L>!e*9Gx&j�S�z�Ʒ�➜k�"���L�� ����Xq�CJ�i��8E��1*5��V�@�r�MN�F��2�e�����TX���a(�i� ���l�\���(^8���"t>��G"���$S��p�V�(=7ew��Ի���J�vQxh�$+��������N�����Y�G���t��<���l�(�������w^��^�:�ۻjAo�U*��K��� xt�%�j���g�e*�qAA��W�C<#L��#E��e7�h4��@����W�N��0�`��5߇��� RT�LQ���WvX�^K��"��C%�3ЎߥYPf����a=�#Am.���>lJ�'����<��q��N����b��<q�:	�G�
^?�e희�Sv�R�O��P�t��^f�m��N��-��-�Bm��sNm;��� 6
���qr�����i�PCB��U��Ag����7�..�OΕF�kp���2��x��m��=��m*��~�j��Ed�����@��\^�,%�Gtj�� kM�v�| !2�;���~�"\�&i;?k'VeJ��X����V��_3w�İI���o��:�5M���8��L�~ՔW���]�}���<�|�Q�i���4)����b!Z|��1���.N�G��xZ�g�;��Dz(�_�<h��O�̃�ĕ�a����;a �R��pd10	؋NK��Ǭ��Sр�����R���4)�dO8�e�	��^����W�(��W�Dӧ��B�q��7�[%/C<�`
���PYb8��<�wЏY��,�9�4���X�Ȍ~E+N�P���ex�vm��&C >,���S{����EB�O<a�$� 1����˴\m���������l�M��v���^�+I��KeQ�.������M��x�ώ'|���Q�FK7�
��8ۆ��p�w���UEe�����«b����b�sڸ�� �cܴd�~�C��bR\�^s���	��j�DRo�F���w��@��7��KB�[��`���+��\��l����k������Q��/����)���X����`[�/sR�ȳ,��e�g�3N��G�g}��P"�V��~/�	g��ȸֻ�5Ֆ��������6�m/� ���S~��Z=S�`�n8�]-*R��$�G���1�V9�Ҿ�P
J�&�*���l(W}Po�2�_�hRᑱ�ե
Wp�pq7���aT�JH[�����ݯ�@�V'����K�QW�I�DU�h� QnM��>��|��+��_��棊-$QM}�y?����AZl�Ǳ��(5���ŴK-VSr=�ai�I�J�VJ(}HG�u;�M�"#���פ�
�@-TV��{V?������FJ���/ ��o��i��K����L��^�(v8�]���'��J�VO�0�H�N��L�T�;�M1=]�b�Ǭ��9aW[Up\CW{�˯~b�b1b6��s�!,����P4$6�W�-�hE���Iڕ���v��Ia��o�
�@ �7�y�>1�J���e�Dl���ϙ r��m�̌�N&�c?T�o+�.����T�!T�h�3UK=�N;{:b���0���.�=K*�L4r������}��V�ٌ�؋���"����&͹��mb�&U�'XO�%v�`�����Y�`��^h��081�=H�-��	�/����xb��n2˽WA�PVgw�W:y!��R%M`�!ß��7�3�J��Ri�Y��dSM��=# !]����=�ت�׫���e|e���pM,>�*.�C��S�1�!1�	� �ܞO�N�>��ϕ��
� �J�H8��%��y�D�U9(aa���{7�o��p;��^_���u��]/��{��0��6�h�ۚL�]/Z��&��"8����<�IY���K�8�`[�rn�m�G��-�<���]Kt2\��8Wn����Ky n�,�K�<P�O[96EM�,:��r���w����J5��A'$����3:v��m0���[�^#T��nD:��;%"a�/�C!������? ��@����:y���J@��O�/�]�X�z�f���e�W��5���ʎk�δ��.�;AhCz�B�	���w��oM����E�N��C�,!�MZ���K\-0@�.�!49
��K^�C�&��#������&x�&���h��\�Ͻ,�GЃ���\��E�����iC���$��X�Xߦ|�YfڮYq��vd썎�羜_8��O�Vk8�f�b�c��D�0�"-�~�+NQ]���L�e��O"�F-�񪘑�Xzl �u~����@Ozb��i��N�e��m�#r~���[�?Mq�h�&���wI����\CY�/�c@o���<{�$�n�GW(��5P��|Ԃr�h��Ǟ��(#v/�D�Q�:�u�Vyg�ԿS��{�+���A�"*�c�5��r"\���E���h��Y���E�Pf�e�ΜP�����Z�sҸ=bc%]5�6�ܿe�?/t���l�v�m� Q��tY{�jG�����K�6͠�D��ۺ/���g���L�Mo�����s׶�ݐ�\�3�޴��;��5�X�H���i�9�7@���ZTȓD����H���&��5��	���bZ��p%R.�ڰ~�72��Zk�}ߤ�0�r�v�֡Gp���yb)���2_�mT�D5ȱ��ЮL~f���'����-���E�)���j�LR'�=�0t�zV�����Q�b�A>�"	��(dI�Vc E�W�0����ņ��w�w��d�>~�b��\���f�������sP� @���H�����E�3���;��w]�/Y����U=�'�}�a�kvGN�Rˋ��!���G�Y�lE�ު�\�AK1.�dن#��.C��m��]��:�N�H�F�A5h<�����<�Ծ�k3�^�y.��ܓ9K��ֵ���]�����>* �La�x̾���qĘ�Y[�)�%z.DK�B�lQػ�v���yN�vG!�Zp��ƺa�O�֤n/r)���eG�U4�SY)�����/���	�]?���V���ѫ�$���.I-�� А�����ԥ��_�Y�N�;��q�d}�#u/�1ْ3�C)!ʭ�CU��~�����Eئbӂ��E��������M�M�,>$��7d�A���2��a(�1��"���W;<�|�lCT4S�ݖ�]�����\-�As�`��0��ʀ�09~g	V��6bI�@�C���w�U�$�[��oW�si_�*lt)�b R*�~�ZD���Qa�'�w�]��)���%k�|���c~C~���o<G��w�,`��T�ɄӬ�g��*"��6Eܚx�O��i��Ӂ7OP���fƮ
����)-�m���o1��o}Z}�Ӟ��1Sj���D$�����<�,C��a�B&�q�c��ȍ3�G�˓D`ǯ�>�9�V�i�γM��v����i���ھ��I-�]/T�N� �m�ApiWJ5�Y�Xo�ni�V���g��u�ck���8�4��֞K� ��`��asǎ��3�F�Fӑ�g� o��+��aG����%���$�X�G�W��p���wJ�E+6��y�*, S���<ߨ#��@��h�ۅ
)�����B5�-��-��7Zyf���ʃ���Z-F���!o"yu�������O�Ӂ7f�i_��2��B8ŋ_��,F�`����д��y)Ӎ�|D�k$*�&�gT�P����d̋��Ym�%��C���F�+��;������NҤ�~�;�3������c��G�hÞ�B^+�@B'#^��ĶM������{����qU���Q�z�<�>�2n����d���)7Ht������-�?en�Fx�-6oԾna�6$�b-�ٖ�$���b�rgj�n����f6���6�V���}�k����?�mgٶ���0&�U&(�EV밋Fu6�d�w�y��*���C.�!4\p��̱CF�[xUl���!pd��^���r>2[����9�@ؼ^��}s��T!�!b0j�QDE/���J��\�x���KB�8$�֞ ;��@i�ʔθ���~~/b�R�c�����+�~z\s��1��}��HU�P��!�,gy2}����T������/��S`ߝy[��3pu]
�|v��<C*�,D�ɂ�㞟�\P��y��J�O{&Oy��I
E~r�b�;FP��>	��
R�v�zC��k�S%�~x9~�,��u�4뵒�ٜ*���t��$�����ʿa�� �F�×!�\Ft>a��Z�D?�|?���02��t	=Т ���M��2�f��֗�i��`��M���$�x��q�޻�|g���ɂ��7�OU2��g/������	��Ukb�*(���g�$�M�J�0�jw�.���`�* A���}��4�-=���%�!e�)^�S��p�@�ҁ�Ը!c�&}�pg-��  K�!����ԢIC>�-����!��>���p�
�� �㙲� ���F&�c�[����Kz��-��p�n���9�3=�gp�j1�L�����u�7���r�f�hb���o��Nm|�?����f�屗�u_3��2S�R�W�FW����L5	=T�qh�M�[�]@���пԼ�/s���.�#�Э������#�YØF7�Z�=s���wU#c�$2Eߟ�=t��勚on�������w�Ń���RQhB�Z��_a���!����bd�,�N�C{���5w����/h���:���1`����@�:�;v�g.)�ze'�-r�?�5�_��V�ϣ�,���V,@hW�A9K�������P^l�����$Þ�R��w��A���NW�������e�+����� U����9�Qd��઒�U�:��w�t7C����t����ab[�YLr�ڡ��:��"'�7C숽@U���:���6ǖʘ�w�$��ˀ�SúntUӂ���_��P�FnXj0�Uj��-Ӗdg����,�=��-K�_�G=_�H�ό>�(ߏ��o�Ci�1��Ð�}��l���>�-�Z<���K!P�����L%^=S^O�%�Ǣp@H�wts6׬_F)�d؋��ѓ��I>L&1���r7�����H�t{o����8>��K�^�L���'K��\��}��Ч[$sjI',�n��v��N��Xl���*�G|���T"8����@���Ihs�Mg�A4߷�NiO�8�x�����S�(*'�vr�;0 �-l�*�b����n�ܯy2�K�y�w�v(�v�+�b�t��i�]seϴ6:�����,��H?b��+�\����˹���F��XR�o����=���_H�#����S�!dd.���:��@.���_�9�/���S�$	��xʹ,�vؔ��#%xn�K+�E��)D��jq�qH$)������df�ua�p�Q!���r�-�B����]���`�4��U�c����*��U��_�{�M��d]o�ӆX/H���c����|�P��vo��I'G.`���I+a�O���������c��4$�Z�S�<����".0�z����"��o3��/.��<�qtS#ۿMcQ:��	��Nչ�V�I�ҡ����F�U#����(����?>k����Y���9}-g�I�G��d�����	Z�Yg\[}ao��E���j�L~�"��R�45q	�8���qv-!��п�������K�^*B�������(t��m�NY6��^sru���P@�EY�=����*�f!8{�Zj��q�;SYA�MvA����#K�S�%���T!j�ɗ���!��)c��$�F����D�]8=%):���]���n�EU����͞F���L%4F�k',�x���}N�(�y`��U����N�'_1��~{��)k?0�oT7=�B���+!��	q˺��TĬ/ʈ�u��l�'�E�}D�(*�ϣӃ�VSa���>*�k{"ʑ�՞��wo�o��W����ۻ�Π"ob�.-�s5��-�\��(�|%�et�Ϻ����C� a�n�ʠX�'�ˇ-Ưnt�g��u&�M�1[T�^ZfL"�`���3#�&�Z���z>���å�0��>�H+��.�)��\��(�j�D�G>926��`�]m�n<�eh>Iي�p��6���E�K���L˜����x:���/����/��Ë� ���$�ؓ`[Bfr3���%1X�r���:�][L��Qs����iժGe���H�E����EZ�ة^���S�����P��(�?�,�/$RV��l4�Mɂ+�\��	��
�[��6k5����$�Π�XZ�7�����:��޾�)�*%e���B���|�m�U��!-[��W��t#r#FB/R=6K3�]]�q��O�������?��m�EZ���񸁪�qҁ�f�Sӗ'g�'R��J�����)�����.˧���p^Q@�5'7��Cў��-XW"E���Q���0�,��zJ��&O\b�"2����cA���w�%6+&:��W}m��X@f<B�TURnz�1p�.�_�7��+f����u� ��f��M�3�{T�.������>*�.r�{[�翾ɇYՔ�ِ�{�H����.]�h�Q�I�4��=u���Z=�<4��B�vyW�����7'����ḩ�v����dٿg7Oz#����Y|���h,��[:%*T�T#�����VBx|||v^�����r�ll%ݪ�*釕�p_����^9����i�lRb�S�,-�0�!g%Jo��\��1����wO�#t��"إMb�h�ї�@�6@��W3���c7��0�� Gw߇scI���K��o1m���`oM���ͱ��_u��!��u�H3���v������:���\:8�^S��&c���G���gV6�S}z~6�-B�0�r!�$�;}1�r� ף�3dYP<}�5!tC�����Mk˩�9���#��K�0kj��~��a�(*UH���F���Tq����a�N�=��)=�K�}U�,�P�,R�B�@�D��P��̀_�e�DԱ�l�D<up���y����,S3���3S�+т�0oU�v�</Cq�`w�=�l�i��LZ(��IC�&��)��to��Gd����I����-\xWv�#�7�׌p��84�O����i�w��G$���i��]���"��z��
�*�����;�vs�Kٓ1{��{BC�(c�d��5zr�Fa�z��!$Ѷh���B�=�uݓ�K�P�q�f��+:Q,x�̀j9��1��^6��`��X�)5se�M�蛼�_����5!M�����o�=Hl��ٔGp�@~� M�.2���60�KV��8K����5?I���i wɲ/	m�ϯg�D"�k�V�����'mcyZ�1��;ɳ�*��0�'���C��2���ܿ�]ċt�n��h��[B���O�W���cq�Zyg{T��X���k^��$J��Z �W�����W^5y7Ѻ�S�N�ٝ�]P��9��c5�|n���x�rv%7�'M��
�+B?���5`@�=��=B�b���l��ʞXե���G(��|�[���ۊ����Q�G�R"�r��#4z҂jV�ڰ�ARt���oQ;��#��6PI�3�5l�U>�Q�_��L�X�l˖.Ӣ���M�D�_�E�ːlo!
k��Ֆ�/w��j����u��R��g:�1W}?CT���0ٻ$3�+�o[�ߖ�b�S �������F���C��=�Y;l�Xq�=����\L�r�w�N�v�	tR;mz^���Ľ]�[�ys¡���>-X�I0/+΁km��0f!�i=��H��ͣ����\�P8B=+��ӎ��:�b`�34�ݸ�_�TY#��$X�wG:�%��[1<�z��,�g0yĐ6�ۏT�X���8q��-�i����"H_^�:i����E����9�U�X5��<8=�mƳ���uS�s}d8�їC�Y[[M�� ��y+�"���'fF-.�cl�ׁ�n����( \4��'萆JH�ٺ{&�"8��s��Y
f#�D5�Jĺ6�ct��6�~��
h�[�åo��g��D�-�O|�|z]���C?dS�ioC����a?7��#���A����J!��I����H���3Ctm���M��i3Qg�'�����S��Nϰ6%�.��BU70U�mfwr1�5G�
"2����M2�o��Ӎy�RM#n�ֶ*�w$/��"h+d�}���4�s�μ��no9�!4�3G�����*du �q�H�uą8��8�I�Dǔi��P��j�xs�N�<�\��j�Z�SC��%EĿ�Ee��A{�������6L�5�E�ep#�]�9��7JȱD��qWQ(A�	�V����;��i�|`�C�4=��1g�&���jA����(t�>;�\9�[�#�
��+'���%_(�o�¨m!�S�#S��96� �)�&�7p�Z=^ի��c�f�x{F��m�}�[��A��჈4�ٕ���Fi���z��BW����W��E�}����/N���1tpeǌzB���yD�;�=
1P膘�B�8�����y�Gyd8����= �#Ϳ/.����g�aS�¯����W��o�[�31V>������2N�� `�\mr�:T.� ��BZ^b�������q�C<����6U���m��F�솓z1�5�[܊��B����c+�B%v�q]Rٷ�5���!��� �����/���������N�U ���h�Bec|L/}��̮L��D{��ҵ��R�&�F�b�MF$ChjD��U��k~����F��ӵI#1�(_����?5�",�J)����FI��aXF ���i��'?麌R�����x&V�'	_p��V���dR�Bh\�!Y�]F�V5�␁\ו�T{n}�C��z�BMg��5���KA��Nь�'CU��C����99x��A���a����	�V� �>���qm;�w9��.M�U���ՙI�0׺ϯ�������):4A�$�T��o�WX\+�'���$0�%�f�$�E�M���%�DC�B'�sS��J�21nCxny����ޛ�
A@m�Y�L�	|�t�Le��V� �����g�t���|��B58��<s��(��#s�Md,4�N�0���;:��|�>�D?�:b�7�s��P���`q�?7�/����i�[�ɟ��]���	��z�1ŧ�+�$�¨�WF��Z	o�������G�(����yX>�f�,��N�����B��2��
8g���=<��vݳ����1���k�tb��*}������2��'��#b�sQ��
��.�G�m�����
�7��Н:��8'���F�o_ =���I��Yj}�6����]b�`4�s�L.X��N I޼ =��);D�+��w2ǬX-~����]���������/ҫt:�+CE6$�_�Y�|��fE_85����3/(�x��-Q�/�u/�:;�&��P5U���*���Q$��d.�N��u/�M�F��:�rJx�v�8�x��g�Ђ��9%�Y�(KU��3�W�ZQ����"UْDF���Ϯ��Y�qҎ|�j1y�W���CA/<���P��la4�&�f2'���[l]!)I�#�Œ�s��7pV��L�M�+8~��q4��)�����u]o�r�����Yf�Zҝ* ��]z���J�v����4�K3�v�?��*��g�Ú4�V](���
Y���^+ۥ|3��X��)#��D�wB�#N#M]��_Sm�f`Ӿ?{.���C"�&9P{�Mғ�Sζ�M��|�1���4�Xr�ԫĔ=��/�$����}>�����h��j��8�+�J}7$~)��Uk ���r<H�\��HT4�
) zt�°:�Mp%�����O��Ìf�����Z�z4��f��-�s��g�2ԭwR?|���w�\�^�6N�
���(��%��fbb�l��,k�oU�����by&U�6-o�(3,>wW�GA��=q��č���z2Ƈ_�ko�b�X��(��̷�����Ko �0\���fk	8ӊ��2$�،����lt��\�����i3n��#x	q	�<���^c'��r}<5V���9��
T�x坭lTl��sdq�[$��&���+��ul��:����'��B���V����)���H6�!�����?�Y�;;�pw���c�|�r�����9���*����n!Y��&*�3sQ.�2��a��<�lոB���6��I�w�FP�8p!T�b�������L}b�.-�*/��zl�j$���xOF���9<#����l�����LW��<v�f��pxB?��T׋~�:�$&��6���Rh�GP#-1h�<t���H�s���@Wd���ˍ�fWV,��c�^�誆wa��w5ޘ;>��#\�������e��[f�%29�(�"�dG��n�/羚����0���Օ�Ou��!�)�7���9���ӓ?�Cr�"̕&�r)eg-�8�)��w��Tv�#��*��R�G�����ƭA�B9o��K��dN��NJ���j��n��7뙣��S�|럘�!��@�L�e�ߕF6w�F�jZ�}X#�&��ci�\5��$hb{Z�d<��5���/PG��tПu�7k�@2�����FY�>ђ{��g��W��P�x5'�=xI7P���'�b��m(�
����8sXщ�G�`���ߜ6�#0H��F�U	���P���)��dX�j�겮��`��؏��]Ȧ�`o
���뒪Ygm����+��Zu�B��:��J�Ltyc����$�<�s��iRĄ�Т�nP�P�K��j���X*>�
.�p�\��:x�n�V����� �\c�:/�Z��B�x�B{�p 7��Z�"����~��?����g�Q�Vi������$�p�~�}�sU����q��Bm|��bz �����C����턍 �9�M�Q���8�����n�W�M�%�π�#���f�'�(�tm9����¶}p���F��eB	��v�dW�x��
8@��I!������J#d�F��>�W�j�,��e��t��F͹�1"G3r����N;	���r	
�s���p���`�H�승���4m=.R9S�	�y2��p��v~�P���6����)D�O�E��
�Ӷ�b/�|%#6VP��w6>
iU��;+�����{�8��<?7�4l���5�C��t�]&�q�/Ƌm��_4�^ ���s�P ԁ�H^��RL��+X�nj9�����ɵ��*C��]�p�R�aa�g]�])�Vx��i�E��L8�ۢw�U�X�P,���%��cG�y�zH�Su��5Ĳ�-���H��/M�U��T���X�6���β����u-�D0z�+/Geo�|vi3��&(C���2 ��X��DLtu!,���T&Q�����ܻ��������� �(;���Z��V�(��Q���:gV�4������]خ�ﵬ߁L����Z�O��du�6:¦�mA�c�S��uΜ�j�qlcŹ�y1�(��D�K���O�ǽ<E�GpQdğ1x[������-�Mvv���9�%�f��a�q���vY���i�����=��w	P�6���:a�RZV�Q�kP�W��K�d*	�p�/���#l���7-��f,H��TA΅i�!�.UV6.�^�~#�e(TyG"��R��8��Үtc�̧@9�tC�h�6���A��|��5��
�<�M�����0�|N�uL��s�hƀ�����
6�`��pi�:�T�Mv�W�N�e)�p��e\�5�=����\2��t�E\B�((g�#��K��5�˧R���7�e}E�l�^�⏺�H� Zt�";bq�j:��S��9q0,�u�-��>]�	��ct�M�d�ek	�5@ք;��h�f,���2-�0_V�Sx`�]v5R��Y������ǶNj
j�"��	XJ��C��PrL�	4ob�U/��ϩ�͒�w�۽�+�t�D��kZ^�0=���%g���@ru�Xy��5T��R;b��w����+�I�3I�-�T!ȫ�j��� S��%\��hG����֑�F���͂�U����{N�L1_c?g�D��h!��o�;��dP�>rQQ5$�Ct$�>x�h3�	����s���I�|�'��D�~�Q�ߒ�����4�$T��sV�K��e�}�G�u��AΫ�s�((yJ;ʥ��x� ��+ѥ���)��,Z�[u_�h�x���,���ڬ�ڤ#1��@�s���T�s�xI<�B���J�p�O}1����b�nm�4m")ﻮ~DFI�v	���W\�x)	NY��~oT�� �"��a�}�nE��#��9�W1�NJ-�Mj����<��E�!6�3�lܣ��
-P�.��7u���O6l{�'^���<�x�B\M�%��U�:�嬆x�l�Ú�e�v-���v���=�˺�@ &�-l���A�׼�.1֖!�ui�������|5��@*�� J�-W���]���Rﺶ��Ϛ����Q'���+}&����1b
����n�����ʤ�䍵�oK���?8uOn�9g��)�.���|�r�" Vį��Li�\��p{����SG]?���h�V��8�%Ն^+����������q����_=�~��3W�Qi�Z�T<�p��Y.lQ���;���_k��0���v{z/	�S"ӻ�\�n��y+�wj�O�C	��1����?��#Z-�vRK&+�A]���5�̴�<@{w��SunvX��,IA��ߩ�hh���f�XەTI+������w�kd)�;�5~��G�`���o���3Z%z�,��K4==-=��].P�%S�\y>FO��&�v�+���9
\9�=��d��+��`�%�#1�-uO��d�&���L����%�$�I6f���FJ������W�w��[��#R�L���YN�W���p>��B��u�+M6#�q�w[�/�
�M�Dn��u�x��cu�+&�Z:�<h�㳱9h�%��ƏƔ:Siu���cA�ΑlKZI8C~�F�:���)�6���9K�z�f�1k�����|ˢބ��l[c�&iEt�A4�[l�9���7�����z5� ��~nl(��6Y�`����r��qB{��m�2�W�X�<��G��.���ڏ����}�/䭫]���à�n��M���&�
W��sO�s/��#�H��^|�GQ�?x�w��/��߮���lh��j�{�w#�\�����ޟ�P����;X����Se���V����7%�j���8�4V�w >bC��U�m�]$^Wk��a����۴hι�����7n�7����I6�H c�y�x5-�K��l`��Z�ū8�b�"�4�����ou�s٤�J�|A~�+9�߼1"�Ĺ>�K�0�T�}�+v�i�!Œx��R���3��zQg'�G�ք� -?��#ů�H��3!x����2=�Z��U����}C.�j;�=�; �だ�b���Ŷ!���)�KRO�d�r�+%�7�LC�*�{L�N\���i���:"˻Up��/?�Ey�9���[��6y��9Ϡ��Te�^�-WBl�咉 (T���������d�J__I�� &U��*�BK�cЙ���ǟ�*/e_`4ݩ�lR�������I���H_��i������l@=ig�������o�`a�`rs"�}	�ժ���%�$��A���	�u
�S�
Oj-F|���GNm�����q�	�x���ї�A��$��~��@{?�Id]��Wd>Ϣ>��$�*����ѧD��
�>ʜ�2֤S�C��o��Ē�[P�7	V�-i<T�I�yM"����[�P"/#O��ٰ�r�(��D_�<��&F��k��(n�=���!.U��`�@�`�p��&ޡf����e ��;��-���+Ȝ
���t}�J�;5|���:)	n�%�ػ��a-c�j�h��A��/i��8�(�5���:Ŭ/ď!z
v���pr�=JUUM�y��ZS�2���C�'���0�Հ���]���_�NJ��:�o���emз,'���K��mV��Nڃ�(7	*�u���[�*<P��ǬU�#Qe+�#�(Wڱw�b�2����?MNx/2�7ů�oB1�o㴥�mU�;��K IY?A]'��`5D$ �I�Ƨĝs�h��0��[� �E柫CC:\��4��H�ԟ.va�	���2�
8+%��Km���W4��rp�� �r�T%K���z��ɛ����9Py@�W+�GȀ�Bu�g�����'��]Y��;p�B�Y���lX2��U��6�|T"��S@���t FVd�,��C��1�i�u��K
�j�K.�s6��(7��N���Z�T�%9KnF�0ʆ��4e: �K��C��ŉl��(���ǭRA4~xx2��e
<�$dGR��F��w�sx�i�m
6X/�[b�\��hsg�5�XQ�*4����/����EY�,�7���v�n����	�q	���C���0dȈ���U�cG�����?�%j4���(&�6{��i�0ߓh!襶���Ч�����E�7����6�!��xx�������P�J�T#�~�jHe��=�qx�
�>�K����C���\r�L�2��� [�A��KEM:k/H��lZs�y�u�W��R�Ȅ��L F�W�o'K'JB�=���`���!��*{��Ç��c�fM{
�=�A9�R���.��#�_�A/V˙�h�z��d2:hu��<$3�������[~VS�T�,�ѽo{���[����jA"�>�p�B��W3U2�d�kvK�ů5�u)G0�0�WS�I������}����a逥��y8�FvR�{�>J-Բ�������0r�r�b���G/.�����d�9ƹ�k���(Fpj�n�;��utf�K��'�,:�&u�v�� (!��[[�T�� ���������-q���.T�G.B9�K�v�G��������z�$�H[E./7J�Q���%@e7��gyrȪ��U��fU{��@�$n��ՂA�c<����泺���&����?_���z;t�5�ۢ_�'��EvZGRraT��9�\�n|ۧ<�}�"X��}�¯��H������#/���ʗz����G%�j��vQ/1�NH�wųL���{��c'�"g�wZ��EoP
$G�,�Y�zuAs�D�̛K�\ �B\��En�m�j���$_�5���a�"�G{RK�kQQYI�ԋ/��^��DZ�v*��a�W�
H���KC5z��کęi�]U[9 $�gDV�*��
֫b��)�-��N��:�b|8�灝�6�7g̹z5	߀tYh��
�Qm���Ug�=�e�YZ�kU��U1m��7tъF�%�'{����tne�-����b�������X޸FA�n��ju���ZB�����aIV�_�Q%�X�tUo��2r'����8}Ÿ�A�\{C�|5���D�'5y�u�7�kW�b
�ֻ~�芃j�,�:����� u��}�5�������_�UӸ�<7}62S����/?�r�ޟ�u@6���V�b�����5������xV�4nW���(DÕ�V��\#�������6�m�(ǀi�JĈ�9���$�[\���]Y(�y�b֌��@��rrN_�R5AnG�Et�$��"Yl�v��Y'�
xic���e᯷�s���j�7 jf�����@e�ۿ>	�G-5��ZЙ<���'xڛ����Z>'�k:wH��l4+������ЮD@z���\yR�`�11|O�Ƞ��&�^
5��Yf`T�5r*���ELF҈�yri	��x�s�����zk���g?�KI�~���h�`L���-L6  I	Y-f�����W�y���,z���74�k
?I����?*R��.&؁D��J!L����;b�4osV��&�1��5��
���1�����yǈ�.��궟u!�.�ѱU�]�ɲ���L�l��L�
L���F�X4�����/)�m9�kf�2���,hU��qi�]Sʅ�ʻ�fS��^iM@���H�:�,���c�]F���Rj�N�J1S~����R����hٖ��7��Q[��]�v��ud�&7lK�����%\W��OY��DI�c��y� �9@����]�����X�s��aDi���S��&jB��I�ӌ5!���^���ٯ��N-=aյ!���S��r$(*9���b���r1sxU/�b��׈3����px%Ѫ�|���:�m�t��Z����e�:�LUф�,�@ke:���JbH�t�į6��h�pjq����,)2���9�Q=w��#�����'���m{c�O�(
�Pߏ��9D}�}ʓ�9�u�e���/�649���{v�'����),���v�Np��Z��;Jk���<�h�r�S�q�Yn�WV/"ʒQK"�l�GכY�?�Қ���n�D�ڬ~��O���ɳT�2(Y ���LI����]��A���W,���t�,�@���W��J� r�ie#�TNv=�.m����Ds�����3�Uʦ��hHsv4kT�k�`��
��`]NSfi--6����� 	�j��-���~]ծ�t�^�enFV���
>$n��y�_�����>g��9�����P9�⢞k*�"R!�0���~�Xv��ɞq:N@˫��b��1V�on�����勹�z<���{ɔttJ���P�u���pA�3�@�O��]Z��6���ڨn��3b�=�"�PA��20 �i[_�\���w���",�r]W�Aыk�e�^UK�[�r��+ӊ8�R��0\葆��	s�v,�#��+���ѯS���%�l\vL�y!�Z���C�q�z�T�jA��tC�T
r���r�'gN,S�����z�2ӯ�� �g��wX����fu�k�aoU�$�BD�)��E$�V@��FI�hfÒ𴂳�/Ff��P���oڥ(�e(��M�?G�?����T�^3Q�����z��K��8��
��z��u�V[G|�%N�%?��*���7�D��Ry��$��б�MwԔ)ݒ��.���?KVQK��˶�����8+P3ĳq-S����6�2A�-�a�Z�yd��˕Lv2+5�E���"�ξʟPl�7s:�C�D�`j�uW����4���hk��&��(_�/���e³��a���D g'��M哿�U-փ6�!��*�v;At�]�}��8�3�� ��f9ҳ�M��;v�KVEs5_Vn�+�M}M��ab�Ay%_�0��M�Cw����C�6I��u�*�������ϖ�8cW:��&`��"�L>Fq�N�����#d��u/�|��D�X/P�1>�Y�k�����梁9�7<8�}O5"��)K,_Q덕�`^�c�ɮ�ή�li�IroưE��O��}L^�O!�7�j�x�o{6.xv��U���%Ujq	e�9W���^7����I�D��C��+IJw!�o����*=A�iͅ�4�����/s�h~E���N/仕�2�d]�:�������>����hp���&�G��������NSC���VI<�E'�����pg.o$v����(�����_4Sq�:i�@⻫�j�j��H�����}����BwX=@z&��6�G�S����)�>�NV:��żֻ|\4	\�5|�����:T,F��h��8O8.R�������������O?$�sV�$*�wee����� 3�oyLs�HJ}l����O{P�>Pt|y$�#�]mI}2�RN\`�7#�c0�L�W������xn,$��n��J6M�`�!�ɿ%)�@�)Ҭ#~����*�; /��*\����~���p_�~:���f�	[q���
/*��V��K�!�
ln��v������<^�6�Z��gP�s6�l�q���0���8J $I�I�7]�.. ��Q��Q_'}D���S��9�B��Ӽ����Z2�jو����W�a�8ɾ���)<:����]⭪��s�����xHB�[����u%�L$���ͅ�8Y�P�|���e�$;Q���Y���Z�	K���3��,�n��(CGn �\�A]�bIQ���m;��oG����<�ź]�X��?�r��Kх���d�Z3y\O�Fƛ4[n�d˷f�g�����ߧ�E=���E.���ս��k���|�b��s&��ud���O�Ԇ�饌Va��ޥ(���K�XI?pa�V�Z�_�G֛:��s�f�8���Ձ|���hPӡn*���R`���})Sx'�ƈb����4���?໻2R6�g'k6����X�2��w�y9��`�Bj���w]iA�&���\��:��u���"�.��5�͌WF�(o�x����l�K(�,�`������	XL�U룈�W1�����r�*��,�.�����J�6�����xL���Vi�ÉW�B���!����)�1q�����:_H.7�>�=��SL���(�B����b��:��$������ew�,��U����j�`Ͽ7��'��k���eK�5l/|w�L����؞��P��_�x���b)c��3|����*��)�CK�I��6�9H"� �,9Y��oI3`�Ƌ�G�Fa �jX8�x����m�hE!����0��;��D�*��� �o;�	����-��<I�ס��Av�����wF��U޾�s�)�F�7�z+�C��$�j��/%뢽>9ŵ��Ҍ��E��+Edꐌ����6�4���-S�ߞH�L��贃wO!����ӵ��w?YiL�H�a��!0��kK;4�'s��XD��`�u_� �[^w�D�����~��`����-[����O���O�)kK?	�����;�<c�|�80�n}G������=��Ȑ���9�H����J��r<� ����#�
�U�0������}W�=��8Ë�AH9���/g)�,�4�s�Rԯ�vZ�Շ/�?��EN��K_q=���f�0$�Wed���.@��b|���/�Yu�盇���n���]�η���7O췕���4a~B���"]��T�f����O����oƐ�<�T��v
�PT��ҶwF��O6s%R҉!�{T��lz_�x����_�g�Y�$^�.��n�����/�-`�\έ�9��i����Z��:2Y^���MZ��s�e��&��z���J��(�?�Aa/Cs�I@T�.���wU�o<��x/��	m'���90���f��D0�{��(���c����r6�bB�iyX�=�z��1�������]��p"Pla���O�� E�OO��&�z����v�@p9&��4�	i��p�B�h ~�2��a����?�w�7W���aK�!��8�j��];�J�ǉ4ʼ�{Z��SV�y,)�L��җ��M�Q�a%����/S$��i���6�џ��w�ͨ4ueO���:�����I)$�c��mI�;$���̵f�#	�'2]*�U(G٦��Z��1e�&\1שU��<zU!�F�� �M�R �+�\���b�E����pGc���A�vԵhߎH�B{�#�H�y(TJç�a�����XyBS3���!�$����nl��~3\���,�L:��6��ءe��`Rw_� �$ܖ�n������9m������	WxY�jF
T;5�z!	"]a�j�D@�TT�&ev�'V��\U�E�+���4.�#�	�zC��șl4 {M�~0v��#���i��S>��f��E:���3��6%�������	�@>#�E�T�QGP�)�N����}C�.9�^�~���{�ݺn���gl�>���H���抧���q���D:��ՀoD+�^L����oh�>�%�i��AW�V,��}XD�I��JܯX��^�Q�sp�9Y{E�Zw5"J*(,1b�?ҙ��!5X,B&��#���<�����b��e.Q.]Wvj�II�0�{�ݝ�}s�.֫E�=�U�-qr^h�O��6�H���MY�����>-��Eil�MU��i�A�A�_ԧ�!��.DS"�������=�i_�k��m�M?���ӊ�Jp`\�.� m���@�b�ө�=K�9X�e0�V��@!	"q-��
�C�7v�&?��?ڴ,�W��/�ȋ�b�ۋ�����'�Rn��e��=P.�,��*�у�o@E�l2C��29���]G���,]�a��U*��*U��h�N<���~)��ۉ$��0��C8�,�bm����P�@^���|��n֭x�In[8�q��+ �?��U:�#m��W_MϠL´���t=�N�-�$���
�P8��%�A��-���t��@n!Z�����Jzv�C���ο��f�Xu��-p�@Hx|��6P���[�y��	?��$7���P�(�
pخa�LQb�K�̰��͘��뺰$L���(�&�E��e�?��A���.��T�'�,1�8,���m��h�xȺ�I�*�;�_��x+m�)����㍩)�4�eF<�*�\�>h��ny�4Š�0���Ɔ<�8-�C��>b�[����lM�|��|~/��mD-�;*�ޡJ����x��r�4��m�Q_�&F����� I�m{��+X���-�����֮)���1�[pu��q���$�?*$�0��Y�޴�O��+kKNNG/3u���C(�~�y�	�-��KGJe`0�v0�I�e�G�1�hm�`1>��'�+ӡ��A
�<{���f��ԁ��2̤t���\���أ4��׽ՠq�ap��]"��� ݲ���u�'��7�|y�a4�҆��r���f�H�;�S��W�S�Yjd�|-�]���BPs��q둓����Z��f l�Ux `�~�p,��*���D�`o[�1������'�R�� �O��}����l4B��
�qa�N@��J(M5��)A�~)zLF8�O����T�Ւ{{��R�)¼�!��ؚ�4`EN�x��ū��.-�ȧy�^r��~?�&�Vf�f˸L���u���	S<���@Hd���"dLKnMaɽ���T.��Δ��J�"�~��k�<DF�1ʬ�&Ǵ0 /C�㞙�^���	#u|��+wP�r98�;]�k�Br��f&���B�"a�4<��I2y�U�$�rO{܅\L��gx�%!� �����l��U�t
R�w�c�z���<�Щ���	���v�jNG����+��l�f���&����N �a�g%>�M��yLp!�')'���s�͞�	t5�	m'�ߙ���',�c�O.�?�n��Gt��Y�n��泔�P�ߎ?ӑ���PzǑ�w>�K�4vGE��e vȞ7h����:tM�����.à#e�EC�ȸ�iG����/����Q濡�ޢV��ߍ\���S�2O�E�{�&�3t�:���f2�:���O�r,~n�$v�M1#�o!v�	�=�����p� 8��$I�>���E�����!�ۍ\�1 	��9��r7��Q����;Kt�[�����2֛(�E�+eWQc���Iಿ��L�t�dі�4?�on`l_���Y{1�h1P�a��f�hܐ�oE�KC])tޠN%\�r�L |چH����F�߲qT[�u$w�-��#vY��M4��u���.�K\�"EG�5D��N_nW��5����~�|�ޫ�	>�xPK�X"���!��3��� ����l�o(d�X�Ji���R���j��'�H��l9Fk���E���&�b�7���O���x��
z]`����N^w
%����{Kl�/�rL�S:�t�x`9�� ��O�L������>^6=fq�j'X�:�ZDѭ5�$5!�=��-��t���*�QěXB�������M+,�I��aE
!�$
6���]�@�b��h����j��溘�)|�������]ȼ{ZruԊ?���j@+J�u�T4M�5��R�>�A�=�2���EB�т3�	s`�����L�?K���Du���W�V����r}> �ETO@W�Dv���#e[�TwZs��@��(��rt��<�X��Cr0��Jx!*��V�D:�x��f��ͨ�������EQk�;���Q���6�"�H����(s�n����l�ls��-����}��l�C���/C)c��`E�ɟt��=�� �dnqV��m�R�Jyu�ˋKKy4.�dC���UBZ�y1�F����+t����0�i�\iĞ�a>�? �%+=�=a\5"bj�rh+�)kF���٬aܹRi��)�HI�|O���}����`�(7Z���\6mݵh�0Jv�u��7�]>��9��{;�DE����y��\)�j�Yɓ8�x,V �n^w��H��X^���@�� g�8O�`C����턔٥�zr��r�+�4�ܾ/��J.40���f{Q��9m����}�q�$� �i��S�tŝK�Z���N�
0P�ܝ�U��p���~�/��ͰMK�xh�ʢ܅	����نW��)��jRV�Rds�#i��An�9FG�n)��{��STkw���:�Q,�̑L�q�lX�I��bu�}�wi;�ǅ%��V{8��U<B�Q���}��,s9
G�����C�xoM���ؙ��z�e�o/��8L8n��g�:��{tE��A2`C��{MqU<�o�'�U,i|����I�$�vc��/Ed��렝L�����wG�JZm�a�����(ʭ3�`TnU���>�9Ǳ��[,� k�pǢ}���`�����_��4J�����+͜���YYj-�|���O��ˉ �v��G��dy�u�!�M�eݏ��"�Ux0>��Ǖ��^��e³����U}��UGE�����-�	/��M��f��=�Rd\�R���2f/qn;��Z&�����W��c���HN�)ݝ�������zjt�r�Y�S^;�Ӡ*���</��i�L�E�f��%c���~l���ThO��R�}@���=�o���za�u�Hɛ�H�(�|ϵi�&�UŅg�Pi�]���u�z����Rj�-����ƴ��~��Tc��n���}��!?6
RV}�!��y��F�t�m�JOC��r�4b��$Y�ph��~�Ї�j��o��1z���>4�W�u.d�'����Z�ej�T��A�ǌ�(�"Oc`ɺ�$�S�]��r�ס�9�d���ϼ���}w)�ǿ�'��w���qz<�Vu�N"��Bj��2�o�F�:*��olAt5拷��rV�D������^-�5YA��cüCMډ��ңM��l�c�q�����n�8`�`n��hgG]�������vB[ʙI=�W�����{�!1?q��d�+��d+=�����1����5G���Bl+6>Yύ�7� #G�U�>.̬5ȍS�ZI-�)�eo��Ā���~P�x���>�h���jxN�z�!��k�z_ߊ)���-�Sτ��a;�oP����WFG,m�e�sd��`������_�^��]	,C�}�ɕi��q�}�h6�g�i׏+�c���m���_���8� �9O���.B�wΈ�k�Y&
@%���@V���{�R��>�C�a��X�	�S=�\1K�7W0�Fa��8�w￨K���U�E��p��� d�\gj?�������@fw�^�sLI~�Fy�(����m���i˶[�Nf6u4H��?(��h}I����w7����^�R�3�������7z�B��Z�+���]{�w�~t|f$��{�˓/+���7�x�;��ln;�6u��׺��ҤJ��R��YCF�DǙB��XR5�"@c��a�&�`+Dh(���'��np��{����� �'zȏ� �=�~o�F���hz��Ys۩>Lw���@{���齄S�����Xo���L+�<È��.8;wk|>��^��n,�k~�s�=�� ��t���z�Y	�Y �ʑ��4i!��J�n�w���剆�Yj��f�zg�2��E�?Fq=���袃�Rײk��ҷ��l�dH�D��W����^T1��ߜz�<���~ci$v���R�i1�|�|��6F�VQ5��A/6*OVy@z-���Kx�B�4]b������_Y���r鍂Wn�վ��	|�s�n?PX���B�Xt����"��6n��f2B��Xk�}�h��Y�);Ek�\N�"���-}-�4|hb�Q�*�+FS6�;���gX�w��08-�AD+��tsZ�}�腐Mz&�ځ �@�"!'���\�I Y�Im#�aE�����&�����=T����6)�[���'�܎̳�/ِ��ᄩقǫR�B���[���?�WsF>e)���g	w)L��w <1o�,�F��&v��$�����⟐�j��D+��r����(8N�(�a+����M��̩�k�h���>���8 m��I��i� ��pZ)�7�5R��fK˴߆�x.��\�w-I����2D��<O��,'���&j���*M�E��, %���58��>��PF�*R� <`}&�YR-�ʿuʁ�먍�r�Ѫ�O�ld�2J�oy}p�Ù��@����$#l�A���v��F?^���.��|��9��P�����N#�m2`���FR���l�r�J3��V,�Svg>�29��+i�2=׺PD�^jyx閩���v*;��s3i:��JuK�LH��{�,q�*3����+�����ƪ�?�R^
����/,b�Ů��4��eSwcC���\�j��Xɳ�\n
A�^Xf�ׇ�v�6)>�_��=B݀4��n�v}��|��f��hy��Q2Ⱥܬ(^�X@e�����B%���l����B
�aG�
*���?$.M��Xk��璦ֹ�*|���q�w�4�,eã���XdzH��w�Wh�4��o��\���zDM|�U���3�œba���V�q-�~�6�8RT��Ko4����h?^@�
x({���`[���d�P^�����%Ӯ�_;5H�C鮎;z��{>!�ط0F�<
E��凔b &�S! ������?�O��SeI����)S| aP��LW��3��"�Hܤ4���3$�o��,�t� ����v<���IP��	]Jtiĸz��蔞 'Ǫ���W��m�����ef����I�G�'r��\0J؅zd��hߦ�򊐓	�ɟ,m�kc��Y?�߮����v�����Y;Zs�+��8=Z�۞�(,��T�ۗD5�f�4�d��(�����I��w��
�>4�������-��X��[:��/��Y�"��Ur&l�Ժ1:�T�j�V����N�@���_-��X?��/�rǨMZȊ���ul5Y�xٔ���G� �ˢ��f�0S���f����ˇIc�SA��y�&�K�)m�C�b^|����%��K��X��I�0�.I�u���*��6T��gܻ����ܿ��=員76p�8���<���Z�cC���}K����|	�K	�wgږ���Mwd,�|���گ��3ÕoJhǠ):2����UY�d�����3k	�r�Pq2{}�s�ǔb���o���ܑ��<�r�b�E�	�>u*����n�����s��/�
��)��ɵ�����]ֶ/?ik��7�Ӄ�ǖ��=?o��O,�L��h�N�K�))��7<��l�xV|ǁC ��ɅP@_N���4тW'�$�yc��/]����z�?��?�.;�,�/�YJ*�#��S?ܛ���[u�ޣ.�y��]+�7�0.G�{��A��[Yt�f�8ne��ѩtE�:|�G�A�My�U������ǖ$ݺ�m�e��b������Tӑ���!^^iogR�kg1E�8�Ҟ}�F!�&�H!�'��#+���4�h�>x2u�O�}%���g��.��s~�~I�8yTN�Č[��4w�g�4sfL���(�uw?�-d��G�OW���?Q�?8�4ؐ.��3f�Kъ5�V��
@��3]��q,�9�t9ۉ�sդ��2�΁�3l��ȋ��4�BY��m����1i1���N����������q�O<#���54�����x�X5�s�\����w3�͌�����D��K8&�확˜�&9��Ű
����po!$�An5��h�<�pa��QP-񟐥���\3�'�G�0��gs���y�<W���B���7��g!�2�G�Wt�	2S�9�5C�}��G�N/�9��$@�.l�Am�F�� �P���@fv��$ �a'Y5U�ױ���g )�0�/���3���N�Ԟ�.I��s�c&���Wkh�A�K��AV!b\ͨ$�طS�별6m����Q�����������΄ �$�9��q���h��;`�{�,��D����8+Z�ӈ�S�kȿhƪ���1�7�"Xbl�"J//��9������_�G���V:ʸ�(ц�dT��ͷ�ZT@��}^,�us"7Q s!F��/�[ϖ�E�S�Ϭsx�Y���q�I��!���F㏰@��w	�5��=eEyFQ�S/0��_��~֬�[�V��AI���GN�)V^Ɲ�XhQB��`B2�ޗ�\��/���A9��0����∞|��ދ��:)��1W�Q"���_M�F�\#�W[NGU��kD�=����_�z�Ǝ��g��!J�ߜX�0{�QD��9ǥ@; ���K:�hPn��aG�1@�IB���d~��7:|�Hԥ��~�pܿQ�uzx���x� ��R�8��oxs�B󻸒�_���>-�Nc�gG�t�Ć:G>3!X���5F�_yJq���G�_��+pR���Ub����q(�|�r��B��DCZg����m��[P55��u��\_8o�����W�/]W�iI��q���;ad�����#�Hq�]�XR�Ɉѯ':�lj=ȝ�k�y�b�o�v�����~�x���9Q�A�''�X�^�EΑP6��	>��c���h���d/�e�� K��%�/'�sG��w��j�G�;r���e].aXҿ���|�='���cb��e(�or9ڇѧ��r2�u: ���ƾb�e�	4����}T�����57B����,�mV�����+'��'�?Zמf*�脜�<[3�e�#�4�4�Y���0���vԻ>g��Hr���Y��ʼჶ	�2���1�)�aI�IQ���� Ǥ$`b�ja��M�tU)��A��<`{r�c�;n���~܄7�����(wg\��`̰>u@K�Ґ����ʌ�WL8bn���UE��/�g�i����7b�e0��mT����A�U�h�x�E{�.�ny�ٜ�����	E���m�����e�o��N�WT4����a�@i�k��L-Ͱ;�`��Ͽ(���ysUvU��nR"��i�\H���epv6���LN��������LY�G���Y��������/,�)�-D�����]������0��(��8�_8.tx{�{��4��K�7�8[���,{�8��XF��'�խ�W9���b;z������S��`{�9� �Gp4�n�~r��P`����n���稗�_�լ,�#����\:��Ѹ�_gJ�q��9 �������}����FL�'���<�11ɉL�*?v=��M�f���*�%��:��!�u�\~FY�J���Q5wDMy2��Ǳl�%��3-�{K�,�ɰ�P�t� pb<aU1Pݪ!�v�p��_�^�ہ�����E<�G~o��90{r#g$.+6��.��㬨URc<4�
��I������g�{I�C���̒E���y��ޮ�E��p�t<X�r;|M�{�1��zTv������!��?m���q�^CZo]*{��%@��у c�I2$�̕Xfk7�H��H�1�U��?��Jܦ�U"���14� �QJ��k���k@�#uw���]�>�����|��Z�����&��o�6U,o>f�Y��G�[i���%�:���≆͸% �z�V�$ݚݤ62M�	�:}�x߶9
g]��`�%�)���v�9����wm���^�y4��:�*)�8�q-f�>ڙg�����Bax�+�ꐁ+zb�q��ԧ�'z\�<����M
�Vob�A��{�(n���&�N�>���q[�y7�n@.p�HS
�\��������{�T5=�j��zp�,ĭ�|�	�:�#id�	=D� ���X�N�~-1�'�wB�J��ʔ��SE��h-�ZD��	�����)sVH¬43��V�0ҷq����n�y\*'�竟�b�Ua�{;�����ɓ�9��MGD�ޠ��v"�p��_,��`��3�"� |(
�+����x�l�{^$=��\�jM��꿦�x�k�^�Ŗ	�aAκ��Dҕ�*�*�Ҁ�����d�xЯ@V��������Dh��pEG�`�
.@�74���.א���+��m�ө@�ɸ>RΡQٛ���� ��!�{
�tײ2��hm�%m<�AVB���_i�`�8�q�.����|@T[���}��o�+K�=��6�sc���G�]����3��5Ż�\���qf{���2Թ�R�zDd��:�ݲ+Z�֚=�\J�G(�����$,-��;��)��b	8�+n3
�Ѥ��X�&�z���ӄ�p�,)�Y��u������m�@]�ܾ �O���cZ.SC�1�����r]d��u�<��'m|��Ԁ4���k�׮rV�g֩M��OW]�=�9TD��+'/���ђx�pkW�,�FyZ����$"Ƞ�{�K��Khyñd�D���y�B� v�7�����֛h�ҕs7�ĲD��cƒDX�7���TA5�3���?�^�I_�����)\��3|��fp��- ���
�����19*
�����N��QX����j���֗ Z��A���hS
H�v�K���y��W�b�����]R��[����0�H|���X�i��>(	�;�j�X������m�A�E�����@���A`s��fJ�ĩ��/U�4y���
�m����V��H n�*�c+�؅�{|�W�Gd�u?��'��&�[W����F� �ǥ�T���S�*�)����S�>�x�~��ه�a�[2��A���ݣ�g� �5�#���$���M��s�O�>1	=5?|D��5���rR�a�k��k��"j���ܩ�!xL�!���)�*z�����`���#'���0^x�Y�c�7ޯS����E3�ai���R V�Q��.Od���ȼ���B@'��Xf�E|��s�X���)��.^!��^7��,NU3��|̵�"Q@s�&̸�x��r�}op�q[����!x$�T�d����OӠ5�[u�w5Vp������G׈�4�L:���+��A��\|[f8^�09�;���|��	��-Q���T5I͊��"���$�q$���M������c�b;�]��$�]����,��m��<�ͣ�d�B�Kl���)�VD,A�sB̛�w������G�X�=�;�a��{(T�zH�a7�0f���Nx��64���I����j�b��]ȴ56�y@xװ]� �1c��=�O�p�c�l=ti���cBj��YvT6�)y������5��p�8���Ƥ޵�R_w�6����ZR�9�3�n��چ�L,e���̚ĩl�(@�Y��8[[���z���V-����/T�=���m�ǒ���_l�Ȝ����Z<m<�	��O*h�~u!a����
�~h%$H��6��a��vz?��'	�Q�P%��do��W�\R�Z:`�n)��8�n��qY~)n�c�@╺���k:K3��#uDƅ��=J�`'em�,=�t^�̮">�+.K��:�S-o^{��3m�e!�Ȧ]?8'���������I��>�v�M�6��[��8����9��v����w v�\�4'���p��v��݇,��Z�k�jD����C����M��"��ak���O������MFY=f�'?K������b �m�Q���^����[LO�(�9��lp5gnT���sh)�~�K6:j���߻�(9���hH�$��[\�k[ǆ������W%x�	���N�g�E6���Ӕ��o���[P���d}��!5�%�#�R8�t��2�_'|�L(P;���[�yM������D�j	�����hg�p�W��(ݵ��-�����ޭ��y���>ߕ�wH�$�B�	Zh��H�9��L��be@]��.�=�2ֵ�,����C1M�gT&Z[���D_o�����cr�a�c	�,�2�ԭ�4l@�K���8K�5�p�ښ�Xސa��/XIV�rʲ҅�/c�AС���!\xwA/�t7�80Z�Oɜ��!E�	�;��𶵐7�3����F8�C�3��Wf�`i�Ku&������U�HX��eյ������P[wp��:*��n�NU)~bd`7٣�sP�2Q��A�����;7&�Ot�}�Q&� Mv6���@���-�$�8��b5`���j�����=$:/a�*�%�t��z��ڡ�Qt>g����.��x��9	B�[�bsw����Ԟއ��٦��Q �z�kg�A����3ԧ3cKWﹼw�����n�Ϋ�_N���f��]�pX���4��dԀa�O!�6�sux��3<`q��i�j�-�YѨ�YU�����
^e̿¨����\#���G����N��>��� '�yDD\����M҆��li��}��ξ.)R7������]���k��J���'^2`�r+� �q�粧�]��f�7��<��*��sn��3�&CX@;k�����*B���}`�Ie灨�A����� �05�<�&fR�T�Na��!E�2��<��0�,ִ��:)����C���%�Gʝ[V�

Q��I�tU��h	�L��*���>�0&��7�_O�s��Q�����2��z�����F�W1�����5H�6kY/@C���� .�lN��A��ĸ�Kd8�~�]�۝�/�o��{E�.P�T�fV���(v�J�l�q�������`�n�tS�e��*'�t��̷Ɯ+~���܁���ʟ���k�>#����} G��P�g�%fhR	�]-��^�*�!I7�,[0��r������fެFt�$z�kŒ�~����@�ۼcW��tQ�P� ]a�y�b!�)��Z�U��x���P��[��4;���Q�(�
-C�@��:eQ8^��D
��]��@Q4�Y"�G�nX}��u���D0<���p�]IE������Cz#Я�h%��y0�"L �5`�-�;�u�0���G�Mv��t���rv���*a�J
��Bl��Rp���/来���>	��o.��#��.I΃����xM� �}�����ѮQTnyw��bi���#i�x=�>�u�|�Q��Kd|��h�@��������E����j[F����H`�~�OS`N��l��s��@�\Rm��X�߶�g�X��$)le[T���JV ���۵�{��[�f�Z��P.��K����6~f��*l� ">���)me��: ����V8��r$�(�V�|n�"0����2���5�Д�K�.�-�.db2�^��&�6���%�ۑ��Cx�ҙ@�&3�[�mMl�%FMJ�@c���:��
�r���
ӂ&�S��OR��iYu�T1���{|���2���_���<�'�B뭍��`�@3��Fߑ����KW��Q��a\�>�[�ߊ~5CS�D��sT�p��ve��{݋e@�_M���DY�FRd+��׮4u��B$��GrNSm��n�[�s+�Vm�f$�0��L�g�pZ*=nU�����+�~���AA����u�BrP�Ya062��A��g*��{��|F>g�6	�_�ևT�9��h�o�����]R�yaHm��x�D��R��F��-mL��A�����$P���x�}�b��������!�8=��[�w��\m��#�-�n�<�G�Eq'�A���Ttwڞ	�D�Z�օv}_���D���|v�9�٤�V���)�v�@~p��U��Ӡ�n�����hׄ�@Q9\R0�(��i�&������-���l�<P4�Y���'3g)�xތ�陯�#ehgn'�q�I
�mܚ_���4�I�ZI�A�m�);>oۯ�]	�Þ[4�ZWk4�l�9X��n]X�Ǳvo��2x�1����=��no����J���Cɤ��;ݾ��C�Fi1�Ļ�e>���茷2؊��-�yB݀A��->h�w<v����?B�V��mӷ|UP)��ˌM�+R����OLC�3�8��H �⠑2�K�l���PK$p�d
�b�:j�A�v�{����C���ͳі�!�ݽ�\P�)��-MN���M}v|]U/����+��$�	'*�(����wn��n/������<h�Ȣ�mT��[��l35�&v��Ḩ�'6f.�Q�uQd9�a����+E��c�~�W)~yN�I��^��9�U�Ry_}�����A��3�s��G��Y`�<<����L��S��꾩�8��.��E\�ɀ����$��?���#a�sY�ܙ�b;�lQ�A�N^�	YH��݂~��|�P��I,j "�:� f%�L���bX!�Em̭���%C",��x<�P:��8[��f��`F���7�Sn2#�3�t��'m�)��6�`�׺@z�%�c��z�d!n@�RY��زX YpRģ�b��Q�y�I�8g����Je��DR�����c�A��G��&\ȱb%�J��g��'��$�Kga^����8��������bΖ��cvϱ��}���a m�lU����N�wR����1;i*�f������y�!��A�X�}٢7��3�p6�k4��K��k�O�bC���h��c��O.�Q��햍�ņ�v
4_������d���v��PX��F,k`�����jd���yHo��A��� �et���T`�+�Z���̗us2�-I��
u'�ü�Iњ��E�.{�Z`xO�P_V;�3�UW�ؗx��Uf�V�9@H�V����ɮ�1U:2|}K:� ���E�a����n�ڰ�de�����#��M��d��|��yC�9 k��H4n!2�����>?k
1��vk �$��Nތ�Uy�驦��Zi��aì_��}P�=�PU�2�I���x3��k`m{_z�Q�Z̜�u���o������B���\(�،��.�(l��>&+�^a&�P�	㴦i��dϿ �@$���$q@�1���s`�p`ۭYF��?!�$�d���ܑ@��w�X��U�h��Ӛ׳�9����d�2��v(#�ԙnd)%�bO.��Q=�k�oF�`��ǌ/�_R'c9�A0x����k?����[N�_�QҖ���%F� ��M�C8�u_�3�d���#_�V��aEQ�C��</������U��)�:x)��:�V�`氵	�U�����+Lϼ��C�d�eĞ�d���>�����ڦ�Wd���;B���i�:�Y�?{�,v��Vz�����ϣ�~ʑ0���׻�xtpS���\u� E�������#������ǃf���M1���B�7�ߨ��>�2�2ӕA��n"<���Wd�-?1���O�حR�t����z��9#&�"��@��:]�Á2��4�w<�Z��c�0��s?��(=����gW�ͷ����^�#��f>☘�Ҿ:�>R�a�Á����(���˟����TY#WZ5�2Ne͊��D�i�;�U��SBh��k����@_dB5���]\���ʡ�j֭w��%�:�u�L ����)�x/�ⱣZ�q�q:��8�����d��z���9�{�rC�7���B��&#��!4�"�Uĕ�P��ϫ��)�J])�vSy
�8�Ӗ�+9��n���<w�U?h�K��y������v���i�:#ԧ��hl�wOF�>��/EU��1��Iũ��9�0|�Y��82c�7����:���4���l��᪊Q��)��X�Ww��e�<'ܘ�
��{ĳ䡱�"��.st�r�`ăR�u��$~�;�u{K{cj�v����W� +�#��ɯ��e�,j[F�]��J����O�}�%<
oa�f�kഔ����۱~���M�j�AmAUU�Ν���F�\Ti�#��X�� ������c�G��;�؀yS�~�mv><��?e�Ro����;K��KH���hY��k���Gii�Y���>+:\��Ů�
4����x�#͠|���d5ú )f9F�*Ǝ��ba3�qݴH*�f�o�h�S����=�C#�<��p!�҅�s�Q����ӂK=7�)�d#<�:���%�*�(�y�P���hc���ߵƿ�]�@��؆����VB棍�ónԇf�vZr��7f)��?��-f���qu��C��W��X�t����;�VgNnuN<�	�p��c��Q7��)��sÌ'��WJ� ��O�]�qcl�wz��4��m��� �d$�j���x��D�Ll��>T]Ttm��t�:�Ņ/%��|"�؄��Ts�~���_���'P�t�5Q��[�rL�A��
�FO�k#���_F<9��bB��
U��)���a��T�D
��t'�]j�W-�L��H� �nL 6 ���N�:�݌�9�9�i`���Pe����#�n�K${����U�E�Ȏ�\ِfԺ��������S~\`Llkf��^g��0X?^���׍d��8�&ʏTŐ4�/�Sw׍|�Kw�g�$���[�G�D�������@�"�2t�i�x�*c��AuTwPx�CnTַ:L����M��=~6���1�Z��)oj�� y��{����g�8L�i@%!H��g����F��*oq\��t��^���s/�"���
��6H;�OOQy��L���wCa�mj"�n��gX�p:��}\y���xd0�R�_�2�O\����0	�Q��~Y��4��r�:�5�H⓱�k

QM��-�����s�ή��(/��T����mx9���=���uv�n[.�F|�6�����T����=U:��� ����Z.�[�W���C,����o�6�h�,�Q�U�M@Y)�AXr<�G�,��IH��6�ؤ����df`�9�������bv�>}�7s��#�E'�)����>Ք'����:�$���CM��Z���#;(�Ӗ$ou~�J��I�Q��mI1,5=:��_=����%���=/a���p�j'��̓I���F4}WnׅP�?� �f
�%�dT��-�J�D��&�N❡�:TU� ����P�-�l��Yhۉ)�SVe�" A^A5Cx���L�'iY���][U�h?�t�ET�5�n����M���×�p%zjZ�|���M�]�t���m�,�)�ྃ�)^��P�{����|�=��\��)���.��k�f���&��쾣�r6�=�u�O-���1�ȹE��SM�ΰ�hI�;y7�k�$[��T�}��F,�G:\�R~�X������;z�ԟ��8xmf�1�w����6~�g;���mIX�.^I�;���D����O�y�E��=�4����c��f���jqt��g�Jr��^�2����j��0|�[��W�S��J��G�	��3�~��N�$�������>��
�qW-�a>ɓ�SD<Wc�
Q�VC��ٵ���B��uF/��h��Ò��}�:U�m]m�?bߥ��6P5v�EP|��~�(���V���"��$�CG1X��i�<�`�`6ȧT���־;�/��VdmRF���x/n�ӜB����>Tu��_����`}y�|�����z5~���p:t^��j�X�׌��0Wo��jΜ޷h
�1��	��&%^�w���<N|������;)@���կ��y���C+�C�T(�WwJ�,��)(�V<��ܝ`�E�%�G��%�(F+6�����B�4�������B�<�a�~�7߽����p�/d.�t���:h���7�E
��V �2F-�q�O��kL���[���w��K���L�'T�6QM8�jD�=,W�|�G>�h��#�m/�=xN���?㫼Fo��%�]���	c>�8qn8vy�yM�\�Uۡ�҉��5��F%_�^"IW��M�جt�S:�a���F����Ʉ�J܆�ы����L�:�?��!4"';|V��0�g(��i�"��g˰6���|̊��?��������I��B���s�~��[���6�Y�D[냜_��t��Cu�3Bq#��kM�6T_�Y�=:�˗���_�Id�eE`�z��K�A�u��㕋�F�2e]��+#vQ�������P�ғ�����W���cnH�0��.�����*\M�جJJ`���(d�U�+��j�/��3�^�'y�@�AKؔ��Yb��Oҋ��F�1��\���u:��E�>�����i�,_d�}P��J��]�8����N��Y�ZI�4B����u��/^�����4rJK���0���cF�������n͢���q��r�d��kb�o	��U�&�]�1� ����q[ǲ����腊�k���~���v7�����)�����'���3d�f�M���'N�<I�T$�L�(c��k��X*h

�fa��#ä��;�?	������V6���ͬi��Β����;��2������IYE�m0Q�݆�/�V@ڱIYV;��ʔ�s���?��3��|�
�l=|�y�
�̜;l'�\V�q��[��0�(n\��6P�$~i���i ��ށ��ʫY�F�����AO�ezN��߶��HN��d��US��y�n�@�ƆZ�(�RwW��δ%e�[����=�Y���p?̮����F�����x� ��3��FKu;ϼ���b-����w&��''�2�5;9|rH�Kn�!���3KO�S`Z!�ju�c��L��"���a�Q7���=tjh�� �k��O(!ϭ��ܰ��}_��_x�B	�X6�r�&<q5)F0�n`lAy�ׅ�c������C��*g�����+�5ъ�{��c^�<��p�n�1�M����V-�<�B�7a���&C���{�)�4Ϣ�o�>r���(�~��U~�X{t	��y��.$mŮF�v����O¢�:5[�4r��垖I22�x�|n�KI@R�Oua�@�xY�H�;>*Q��ʋ��Y���I}�μ�������~��*3��x�r���0f#O.ߚ��zᶞqۦ���<��
4�����%�>M~��z*��8���2����:'�cc�
�RT�=*���U�ϊK��\�;׽I}���/I5�s��'!ycz��K�)�.��
cN٭�؃������B��d�B�0�?�mNH�8M q���dR�J~
	1��05�Y|}%j�����9�I�|R��y�;�{�����aW@�Z_�=
g�u���-(��a��R����b���?�a��Y�j|m�5�ͤ�Vd������<J=�U#>�!��|�;�/��3S1��'v��%џ�*�R�D;�b���Ô�t��`��g*��@�Nx� Q��̀&Ũ� �|E�~�3݂�I���r��9�w�;����V��̄�c�Uz��r�6#�<GW�>3.@�fp����"�[b�w����f[�F�+U�-/Mc	^` ��kZx=z�Z7j��������LŖ�Fn��k8��O�P��s�Y4(hx]���{l@(�ge��κ�7Rw��7����$Y-y��L�*�:�	���o$h84���E˃�m郳ci��a��ʷ�c$ܰ����UΙ��mϚms2��7�}��x4�����p���������<D��.��� �+CJ�v{�5����im1��s��j˿�ה�;:7�<���O�S�	�sB����[M:�����fX�-���4|���os&�z�GYD�����R�	��Ρ3��:0u�p책�_I��,���FF�q���x(�?EM9���P���=�܍��	i�\���-�%nף�p�etJ�J4�q�%	\Tu��P�7��v�z�[��P4�K��H�DGq�pQ�]b/- }?�F�]�Y��?�]��8^�)���N����#�Z2�5�Jy����2MTvrU�xCM�� :����������qĺ�\������%�?� ��"��=���;l��|>q_�Ʋ�˩ǉ��V�I����฻��>��BQSU�Q52>�;�'yB�>c�ɂ����.L���k�01��;��E�� Ğ�~�Vod�J�XK*'�f��oc���>x.j���`f������/��6�\�V�%�B��[8�}�v��o�	q��֋]���a�	�Й9o?�ۿ�G�[#w��˳�Ć�ei6NVX�[�x�}���tD<�e�)�uS�{ '5� ���=���q�,���f1�I�A���[�x$�����g�ŐP�so��s���������]�ӵ�LJnw5������ӝI��k*�DN0@��aT@�Ԛ�a�0'R���g��W�*�/��"*�F�J�@��� ���Y���XK��_+�S��Zۡm� P����%
�����/���hC�9x]�z!̧5�J!)^��p�`-a�.&�8�YX��P�"u;�uT��YUhM���"w,�L�su?c[���E�U�����/�G>�ryRYQ��{�6�W�����M�y�J����4�S���)f߸����a�)���
��D�~Dl6V�mB�i��"�!�ETM�u���,[�0(���ڛ�7��R�����x ��A�@`���蘍͜Զ3m��nd�[ �����hfx()JA��X�O�G߇�l���z���R�Bif�Z00���"eH���M�m�ia��*���i�a�.��2�!Z�Ҙ��~��|x���07]�"�O��z��,pU�R?�ʹ��D{d�,�)���LBFNS��bo����n4��˼q-ޡ��N�*;�~߉�BI�r���[5�Eh�ȶBHQQ����e��tAn�ť���L�
�MZ� �t FF"b��} �����ʶ�:#���޸<П�����?LC��:�e
l+Q4�c�]b���fE�N�b
A?)���C��L�
?yXD��=t����PX^�!�
~��%p� �b乥���tA8���) 6=
��#y���^����NmS�����+�U��+�D|�*~��X����
qz,ӟ�^qc�g�ШJ���SL$�F�D#��$G�Ge�nƧa�N$� ӹk����g~rr�0V��&4�K�_�s��-x�!�MK������(��>T�hS&���&W�AB,�"h�o��uuG�A��~�D]�+&M0��Β�)S�e8)��<��W	#��Ҥ�/w6��kh�X��*(��I�z��:Q���R ��3�-�lK7Jߵ~�VC�|�wC@�<�ש�<��f��~��z�ų=(����Bq��
�(��4��+�SQ�bDZ�� V	��	�ٴ���H+�a񒋰ZI�!\��	 �\�����f��6ϧ	X��̸b��Z�Ϝ=�r�\X�(��)��ȧ�~"3hB?�}A�����F�g���b�_�q��Wn�,����p�i-�?�Ti�PBx̆��፹>W��mν�9���Ԋ(ֈ�Խ�}�$��W��`�h�8VS����fK(�t����\�- op��Mk���8W���
?��֪�>��$�is�WFcG��<s�>��F�W�֬y�΀5/��M�"Z~�$�[9P����[�Cl�`���	�2j��K���rW�"V�  �>(/%v"%_�Xߟ�2`��a��IO��F�N�扫l�F��D�%�����?�cDM/�"��=��nL4�E�����@�F?�h�VW���^�%Ae��"�u�*Лw�6��T�{�,�n����'m.5�P+E ��&���vv0YHz��/my��(�����D����S�v��Y�?�����&qiq��F��Z�1�!�!�G"�;[T̪P!'*�P�R?=A��� a�"���$���E�b�Q��yP�!֊aI�Þ���V�th]/�)�۴�>T��=�X�6(�(�l��$�	��A0'r(�:�7�W;Yi�*��܆�죃���[���J�)29��O��B ��,rf�O=�f�u9=�@US����"�Z8yO�i�z1W�z��9,�,l@&j�:��+>-�O�Pj�*��Q{�"��[�����M[Y1%�w����Xo��~Q)�'�$fl����ًHu�Ӫ��j�`#��#`�d�^�V����$� huGo��	u��ّzm>c c�xV�X�3������]�ڐa;�ߍ�r�)�q�=C��W�-��EF+1���	a�����"]\ƍN�!,t/~_�]I #�����GD�%<��x���F��m���*�O�u?zѽ���z��<uI�wn�=ڦ��}r�y��1�~�鹘{�gj6��(z��'�N��j U��(]Ž�	�$�('��l֯
Ac���������Ϣ�әI��z�y�3��d2�d0~y�.Fe	�@�k�.+}i�	�О��s�'�D��e��JH P��C���5x<K�`X�(���f�;���㊴��\�7F�C���	�X��<<���Rg�mdY��������K�<�C\ B�D?��)Z�����N�gjAy�j6�1�t�����!������R��?�'n"�<(������O�k��tgQ����)�w$�g�X �	E$r����y��_��#����!�]5�*�����1M_��Us��f�f�?m+4`�t��¢��~.�W	@|i�?E1��Sr7'���3e�3���87��Bw�������qr]����W�o��-�S�Q?K��#:&j]`�����D':�PPI��x��L�s����]~�%�!��̒R;�^ql���K4 ��V0$�-�D�k��.����w����~��Z73z(w�!�Ɲ�|���TA
c�E�6�5�����'1�kG9$�y\���k�����m����{I�x�j�)����^�Z�]
�0��-��i��u���l$<.��g���e�1P.7�x�[V��βH{z�������� $��&UuKA�S�;{��Dƪ����X̬�.g����FPFhܱtA��s��-|;:ꨇ�B`B|ޞ)�gӶ\��0;W`�0�
�9�s[��>z=d*]�?5���A(��k`�G��'FxH�'|}$�VI��0����o���Bxc�on�퀃%��̱}Lm���	ʠ�X �1�Ӄ���_�c�k�׋�����B[���8�����)��N�
�f���Ҥ�P��а��$r1i3z�"삏f~ؤj�:�n���/���X��Q������ZrOK�YΓ��a}��+�g6\s�CBpGh	��#�dP�=.�<rG*���e�	d����YK�;�k�Z�܏����Q&��v�:$�ƹTZAB2����u���*,�֘�k��p��7�$��z�I�i3ѕ�f���!b�A���eaN�{���9F�9�"a޿���1@�8t�][0,��V�����c><�K���w=���9��Ժ�Q�N��M�yDi�,c��BYJF�͵��c��l��Y�^����+6�2f��M�ǂ �O,���f�22�I�"Eih�2��D8�@H�Dկ�q/d�/u���*�3�x��@̓׬SA6�_Jo�+�6*��o��	����-R�4ڗ�b�oҷ�}�|_��@ o��O��p	^"(����T%�bU���۵iV�Y�[`y�~k�E�z.��+Q��Ӭ�K�2�ZqC��gǄ�����٘e��	R>�2��S�{1�'����%�|F봈�,r9A�c��(@=��2����t��2?v��Fk�ʐ�D>@F]b����I15;��,�.]�W͑u��{��3谮��L�_MIp��I�1�q�X���j��fA��@(,�,X���`�����b���2F��I����'���� �]�����1zl�i�C�{
7�h�Z�c�虸�w%44��lD_V��꩷Ek�I�u��*ck=f��[o��e���L����.�XTI�	���>�^|+���%?��J��^�(����?$(+21�<a�%����>��x�w�Rc�y���� ؂EZ$�?U"�GS�1���,M��<����g�O�(�pm���-lRq�sI�&I���9��G�'(���e �y���'t�Q5�=���c�T.�J�a��(7"/["D�W��^-|�Yz��?�ʢ��,�9&�Ph;����V}�Bi�Ff��E'�"�����͚�*4�VM5��Ѩ��ݣ���)��\�sڠ�=j�$���x�zK�0{�'Ik2�=�7~�x�-Yh<D	�	T�i�������DJ��K[$�]8�i;�1=�܇�������3��f�J=��Oʊ�o��v�i|���L��y�%�������r�e!T�F�)|5�Yr<� �1q�o
��m<��K���%�x����딷'�� }@~ny��ώ��]�ΪhX�q�m��p~}W���drpT��<�!8�J����V���tl���Ͼb��Ŭn�87�`tR�`m�����cjr�Ƀ�ˤD!�V]�£���L�O3�� )2�n���Gs�|�{,�����<'�`
�c��&Yk����L�p�)l]Y{��ӘQ[@� �`[�7s�sM4�ml�7?�e�u&p�3�([�yH��Q��~��b���$�s�!r���?kJ/��#h�DkH_���YB/Br�ɝ�]Ü�М3q�DW�b_M��#���^�,Ӿ`*0�� :'8�X��R*w@�=�Vmc��gю�#� ��	T�ߛo���Sl��݉"���=ʌ�n�&Zܐ����G�Zh�iD� ��+ew$W���/鋺jU���V�j�gjR�0��Sg���x�ҡюU~�3��n��ܫ�&QH�Vڻ����`F�y.�w����*D�����u+YX�����݇����+���Ϡ���Tx'~�߼��Ew��}V�6������>����H�l�TyN�-�nZ��"�Qc��vpg�����@q�����;3���3çlHc������|�wK= �r��Fh��\�:}q��V7���R�w��Y6e��IK�Bć����c/v��6"ԩ �y�wA��a��k��[�&!R&��2���k������v~�&X�Ee~�j�@؁�I���䉅#g�Z�mC.�$Zy����J�i��\����_��'�.�M2j��h��Ԍq�X��9�'M@h�O�p�s�|�Q�Ae��&�3mI���	n)oojfZ�r��l��3y<��̦mi��h*q��\)e	8��9w�������y��_�~������~q�-�)�g��Þ�i/g_O�����2�s�I��s��ڶ���h��y��)��sG]�TUo�#���+`Ġmv�w������LQ'�y� �-������|�N�}������#c�U�ԲX����g��!��`��9��9�},�ל�LOpPGA_����2����Y����G`B��� O>��H�U/܃r�>�˗�mO��<�Wf9W�^��<�dM���}4l}�Oy=�x��D��$ɵJ���h}��`%c~�rDe ~"�Ii��x������b�0�%�Q���Fç}�A��	�('�n��G����^��̶�yս���M�Hi�,7٥��[l����c��ᣦ�R'�_���/��ݖ��\���lF���(UPo'�F�븙Tx��}�q)D\���+Cg���uG�t.}Jo6x�X��b�<���Fa��#�*o;��6v/�Fa�1��t_�K5�U��\� ��$P��?p�ٔG�(>Qd$3E���(b̸�V3�"�N���2E��� W�*n˶A��D�=.Y���*�]���̦į��k�La/��Xep��p��4�N+V�j��M'�8��F�7P�r2:��}���>�w��ܥ�Rs���412�3�D��+��u������r����ss���}� 9�Qm8,S�to��!#��N}�u1�_�>�R�8.x���P`[Ξw"	�6�+9�c��Ճޚ�{�E�B�Y������XvD[9uLg�+^��́���0��K��`}8�p��R��@��>
�P%������N�����}|'Q���	��yQ��k8�Q���~X�P�ɩ�H,��#�����%{Wұ��	��P�OTͻ�6he@ZJ���h�W��ܬ���a���6��,���L�������ָ4 ��q��$��Y1��dgj�e�%�G���A�:p�cAF��D��ߡ1�2k��:�E��޻v��M������ǌ�������w�g*#�߿���'��F	���,Ǳ�r�;D����P�
@�;C�$�Q���@�r�u��6A����v��,�(�@�Ⱦ� ����%j{�5uhB~ˏmyEX?�7S%�u�Ppx]�{ZQ� ��K�D����i�)��"l�n�L*)-}��$5Q�~���+��.ՙ����7h�u� �� =���K1/��r�9gO�GQޠ{|�d�x`Ti�"p��44\�ێ��ښ����n�ScXP�o��T@����ڊ�D�d%!+�����7� ��-R���?�!z�S��]T�إ�@e�7 �|���\�����9.�K4�h&�2���2R�~�=��-��[���r��Vϖ,ǡ@ǑO�f���7���Hł�viL�R����L�Zyctf4����`6�0s�7���!l��0-�+����|�/��9�Z��?�BB,��R'*�ŶMXc�D��k��r��E}�`9&�n�QJ��`��Z%0	f	gw�{KP�3�P��fo>"�p�:�|��@O��� ��?�����=_�bҩ.�fQ-5���Cx�x�֞�.R(dN��ڢ�E���ƣҫ���R1������v��J� |�	7�wr޸�AK��P� �嶸�`�2�-��:O�/�Oٽe�b�m�כ�-.';��M=p���=�b9�w9��s��~W0~Q�6H�j[;��2)��6��@��|��!	Zwrf����'��H|/I����[��a��*����
��Y%���d�t2�2���؎��t�3�C����!���| ��Z��99�Fv���T��=ѮY5�6�F��.�C��mT��+f���lUr)[6J����p�����%3p�ֽsS��;�!��`-b�w�ܼ�֙38�h� %����9m}�1��;�m��6�*k��UU e��������ߗ�uK͍k�V�3�~�����?8n�C��c���b��7���8B`T��[��m��ya";Ѫy���C�|�1i�K�ϯ�׼��1�C��_w��,@˚�<_i����<�0�=�qΕ��-e�	��O�,y�
q3p�b��H�r�g)����Pl��n<n�"I�y��F��VX��.OFz�z*�1��_��_�����+8X����e�uS��g ir'J�[�q%�`m��Ak�vڌ9�ߟ�-xX��>r>��az���7ģ����TID�+�]���6�Q�v{ٜ�]�R��)b�X<w���(�rR��d�A��Z���r���\�^Zԏ��plx��@��}������zm�*S.>�):%q�P��<���`�h������I�b+,��m+>�s$��#�LgZ/1ӎ�[��IҊe]Y�Ӿl��(jdem���-�� x�Y��<z����I�}\�A�p� :�m� 7�ӴP�.;�=�
��Y�R�^5�^��3���s�>�՜Yw�m2jN�C�ރ�{ 9N؄w�6G������YҨ�|��e�������c`#A�+ѣ�Ìe�dN U�H��3���G����=�ǃE�ڀ��WV���-z��l�!�m��X�{C{��0��8-��q���S��,�l��Bb�@�5�wMU6�j�#.���v$8 �⑌���g\��"�@p|�e�h�Ǉe�O[��NX7T�"赆�#�(4���J��Io`��T��"č�i�O@࿪N�]c�e&q�ALT���ݠq��0i�v]��ܲC������`�ӤE��(��H�#��II�]F��-���Q���GS�F�� �����EZ�.���̸R�z���`���-��Jg�����4 %����l!@�@"S@�|�i��.4������#��Xp���l���L�l�$��Ae��3���a
DN� �����58��p5��QI�!�E��'����N���G�DA�Ç�Ey6,<O�DЧM����74⑮�v.@�_sj��I\!>�� -�n�n ���b��tI�rS����H IAz��{.�?k�� �&3�*�Qxsj���E��;�w֖��nM~�w�+�Q���#��H{ɭ\9��-/r��{0-���s�S$��tlM�	T����dC̝�~�^X�6Ņ8�����H��D$��|gW>�@h`��]��x���'���xz��$��J��͎c��E��cUK蔲�>�٠T���x�x(�<C��6
���]z�#�I�9���]1�.�����v�cc�v���L'7~`��'���6����8��V�
etǚ�����J�,�*}�9� ���f��<��_�$�k1,*'Q�!'���k�>�֧Fa'7�̈�����>�� ���so�����t�B
q@���ϫS���f=Q�n��k��i�\���oe�lT�/`���i\LԵ��i�fZ�'�^��<{�8_�^cf7�c��g��A ��Mj�����!ߨ��?��sEj�c��F�3[.�M����\�)��(�� Ur�}�u��Em�O�lU��J��} ���+�L�/�D��w865E�yD*m(7Xfhg-Oa��mQ��weZz-%�eu��Ɠ>����k(�@��x�o�����Rj�|7mP2�K(��G��JI�����%�=��|�n��\C��pÃ,���O�]��C4m%��X���c�ս�I5�|#�Ԇ�'��0r�H�ac}E�����Yd\4����0Q�ސT�_lT<8��]�D� &��y^�%.�$ۧC6wJ�H��jo�Gϰ\w����뒼*BV�+�bDT�I��'�2�,��N����ny3$}�s���c=����yz��#�Rt�v4�ż.%�'�]���!�G�^Q������TKu��Mk�X�Pq�'�0s/R�=.���B�0�y���L���g�ꑀ eTJ��;f� T1�Jg���,��\�a1vg=	[rU���ڲ�*w�u���$a�t8E��`ԉW��R��~0������p �Lr�AZ!�19��N��3h�0�KS�0��a�+Z�e�mc0��a	�\��.s}�?��"5fY����Q���}* �_(z����8_ĺ�`�o�v%�p׺{ ���v2����L
2�
�_Ǜ��:)QS}�Zp����ѾNe�2�5��a�.�٢��8����l�o-(�YژQ�V��jd��@
!i������$����B�>}0��n/)��3�5��pq^7��"/8�T�t�Ӏ1.5w�h-�5B�-�����*�Z��sa�G�-z���M*��Ğ��'|������:~�˃���.9u�?����lЀL��Q�Α`[L��[�����SL��5ԫ���6����*���Pgh��o�u���ͩ�=F�j�"�I�,~�"N��"C&u�2���2��瞇9?_Jr�Z��:�I���]:t�nD����Ȁ��/9�&��n!78 �Ar��!�i���p���0�xf���2�0V�Zakj�C�Q �'��.�����L��Z5�;v
�&w�촁�[ȉ�� �T�QV���K ���6h�6�MRCVRK�X.+8޼��no�f�E#b�d{�Nؔ�����un%�nc���;�$V�e�v�-y�G�Ņ���n�G2DgRmB��#c,��x�%�%�3�� E��4T`��(}[O�v��� c�>�P ��f�qo��Һ\�Y����Vo!��I_�|��%5%L�"�'�S'�g_s�$�d8��:c�]uO/�=��U�GtsK)W�.�*���Y.�ʚ�I�Y�;���j�����j�=Ƚ���DyT)���[}���5S7�e��&��#Ќ�n��gZ�e��bYB��f3pa}�U�2�V�̹�p G��Gnt�BD�9�32�9����L��;���;ɬ�,�q"�6�ƾ,����:��?�K F��"Լ���<���5q��#둨��
«R��ܯ��J��a �qkZ�B|��yD9��\l���^f%j��>�sts�(iI����c!�ýO�f��0�N`���MG2gm_]��o_)�2B�&}YmZH�j��yҍ��:�VlDj6p�6��ٛV��w��AL�D�o*Kt��ge�����ya��gV�Z<��{=k��f�p��繌pc���"�� ��{��ۀ+�%/�8N��0�	�y�������u�_��9��{>fHۮh�|h?e����y#d����&~�Y���t֗f��k��B_�a��T�Ć���z�t}�5GO3'r�X �x�[�teY*9��8ߐ�:�O��ځ���*R�9t8p�ji��6�?j�d-C�xs�&���Y�w°�<���wet�����'�\�_Q $X��bL��(�g.��u3�'��@7��7L�tgChw~q$e����8�=V.>�e�hvtNN��+T��U��TM��2�-̢��ڵhs����k9~�rsF⽐Z*��@�n�޾����]fά�����V��nݨ.�H�(wr�Ɇ����[�1�#�D��@*��L�9��G����Q����ն��(��2S�X	^H࿡���^�������vҌd�y�L��{u�p����[3[��q�ً�i6� -��&@��H�Q��zIj O�����]��+�v�%2���'�[�l��;[JF�� Q�糧�-�� �!��В�u}���)+(ݐ㇈�i��-�"�
C�o��x���X���Zm�ڵ��]n�Xl�{y�;�<Ի5�q(�k�;�
�(��Z��7N�?�1���]�X�j~������_	�.׏�A�4H��C���A$�g��$Q����A��E)�?Q�e��cW��Z=��~CLL湪l�ZyT_�iD�uSU��]��������i�.mXs�zӻ��.ey���`Ԣ�q�,��/Lhn�6�����g!=�"���E��4JTD��)���B��|����:{��\>�El�i�����w��ΘC�v�I��>%�D�:�9��a%ֱ�wh��]L�L�hWr�K�3rkv��ŀ,T�����i�v.�K��^��=�?DGL����㈈?ͳ#�e%k�E ��OV�n�
2!]6z	��&�̓�<{�(��v�A\��`b Ƙ��s�'r�|K�ϻ�|�n�O��s�iS#]a�d��m��%LԻ��� ���A��La	DB&��}�,��<hH��_��%QH%������*��gj1��?�f��+�NO�]����7�2T=t�'����`.��Y!�_�P���]�B� ����y�	��{B�z�ɮ������!�/)�+G��%��t��Jh�mK�/D�g�u>A�W~s�b	;�b"^�O�r�F6;Y�r���8��J���&���C߹���Rg���~oAfAB���Z}-ej�.^�?[丆vYѲ5�O�9lt�yp��T�?d�7�Cӻ��@�KJ����W����Ҳ�in��Ert��LaJY�4��.�g��1^����˭�2ޕ ��m<�E��T+�4z ݫ��ǹ=���c��?��I�T�<��f?�/#�Q��>����D��d��\"���


u'[r�j�~-]���x
�d#�M�+������⬏*��඗�εR�7q��$�H�W�����K?5IuGF�W��S��4!gJ�
)�Tl'��5���=T;+MGp2ķ&�ԭ��yuq�����v��5!T���D#����ߗ�(���	�r�w���2��NUhV:��3g����faM��'(�"f�g��5�r�	&��E���	e�A�s�H��9H�#�h�	�9Đ�}Ⱥ�F6�[$,@̔vDd����p�
����]�[�C�),A�xЛF��Bw�Y���b�I!�		��ә�@�X�N��R�4Y���PbyD���a-gXX�O��6+P<ׂ}�HMGj�����Oh����1�g01�_1S�~��W�6F��{BFˡܽ���%~��j0z���ۄ>'���0�)�cy��β��A+�����b����g̴���qwvJ�1x' A\D���h�Ԭ<4������cq=+R�j}��Y�;ŧo�\SOm�b�g�Q�tN�������q&��$O�~fg|�C��@��%�)�-�䮤�$ �hR��}Z�m�lHVԈp�.����W��jb�F��{N�� �[SѕYL�b�&�nh�?
�	U�KI�R���TSb�R��黚������B���~~��1Y���h/h�0��#��E��:#�^=�s��:V��DA�<2�Ҍ�>��\��Ô?6'��W'&�y��GN�#\��R����$m2^�)|a�r�C�ݗ3�O��]�|�|o��T�-n�6�&�0Vߥ�ݢ���4�j!|g�O��"��^�
~�<����ͅo����W£��cT���b��¥C(7 �Ry�c_�"8� ��S��(���?�L�����e<���h���5�HX���ީ\�ƹ0wZ���{ᵤl������x'͟�["�K���Ŏ��6<�q�R�s����Ѵ��k�r��3��ɱ��'���b��-y��Z'Q�Wv$\՞���+�"z��:�`J�U3f۪�ƕ��6%d��Ɣ�g� :�
U�)�R�J�Sk����>q�������Q�����ù���	�'*CGv���iI��)�srm��'q�LZi����ަ�����@V���"b��A��5���"���Fgx���m�|q�Q�9W��B�Ƃ9��d����$��Ba�Q,�R��DOY�$J�DjN����/���W�}�%$�&��þH��2e����י��=#'�U3��(*��ZA\�S�N�VJ$�g͂<����a�!u%&X����.���G?H-�G��>y�vh�X�$�Z��&�m��
�Jl#˰�������q;^x	X� PC��&i+�;��fAiS����_���1W��.�����?(��$���}1&S�5~ʥ�����vC�-"�G�O���ÌH��v����3�+4��8�V��:�A��bCCc{'kLp��P�խʠ�F��%�iQ�A�B�5;��{hs��������y�Hs�{kƞ�ݞo�iL�X�F�j	1ܯ���9	�f�@���l;������*`�YHe7@�r~"&v��0jj82�i/�j
����!ڨS1�4(�v���E�8���&��Jf�����Z)J������1p���ft콍.&�iP#�W�^���u�c0fǍ�w̞��]�'����`DV�u�R@<��ڽ-�I�_zK��h����2�+r���0n�d�k�@�L�^Eu���%+���n�\�9��P_����� �ݵ�}�O-T���bd�Fl���0�e�~E�o<)��03X�/�y72̞&�S�����٦�T�9ⅅE��ۧ+��m�r?��S�uE҆�A�K�����ň8�t�F�jr�m���)�TY�98��^MƵ{����pâe��ZE|�`��	\�ރ����|�7)��/����jN�~����}����a���J|��p�m���T'��ae�����8ԕ�h�Ȗ��ʤ����r_��-����a�ީ�F�`���Zj�D%��������nmY��4s�t�St���@���#|���aЎH��ܛr��D,�;!�,���NǙ9q�=��82��|x!�tT;���=�B��*�!m-�_�;E�1~/�{O�#���a�p�,u��qF�|B~��-A�v��1\v��(�̼$@�">�c8Q���ƾ����o��X,�C4�椕��[I-�s� ����x{�-��K�T&�2W���!��'!�"5�D�ᡮ��C�(�B��Śi��n��7�0�'*
�/y,U��90���M�����z_�������^�6`7�N%E{N�Ă��L[U�IE�% Vz18&
�dB�,���L`������2�R�9]�м�aJ�K8`@?��}2Y�����j����Uu��ѩ"8��:�\��/�ܵN1�_-:�.fq�4�.o����`�P�ߡ��� ��$q����0Zqsg�($�t��p\�c\�v�;�zr[m��+K6\�jW���my(����Z&�nT*�y��mB:�O��Fӫ@}=��=QgK���1�k~��+���j��N����`�|ڡ�·cU$+�?�/��}�m��ڦ�i`G�*����z��I s�wB�	g��3U��cp,����7�8k���yzH
�P^$�h-�H^;7|�{��?�����Zf�W�/��)נ)L�3��%"n����2�~�/W3��}���ٖ�O�^��%-��K���cc�$?�ל	+d�D�Z���]��=$�ɭ�e�]s�f52�g��H��e�����-����Py�C��]�Tq�|�V���Q�v[��cZ��MQu��1:��F��ueb$���UD��.3���`v[[pXn�`Y�CMN!g��8{�������Ȅ�=��I��`8��+:��_}���uڱ@AV*^�K�bo�s���5��Oq�s�m�&6��&����9+�3l�lwDDnDo�)���7Sbx��W���t���ݶ��V���H��M+�Lm�>h}���@���K�}x�! )[�k�wFI4:��r�G��x4uf���B��=i0��Ww��?4�Y�$�ۛ�l!��z;��#�y^�[k�̶h�+#��*@�x=�Dq�ݴ��p�bk�z�«��[�C���8�s�U�Ѡ#(���l������˾�W�MO�}�}8��t�:�@s�˷�U�.��$7u0�z�q`�3��f�P��_�fъ�y�s`5�E��G�ۅ��t��F#/�(*z�`xV�8[�ܝT��`DO�6��f�%�=�F��	��О��������!���~3���F���d�`�;S2���.�(�	_8����Z¿���X��J��\c�L�,Nn(*@��p����ػ?-l��xd�\�ߜJ�=��z���j8N��0�p��&�yH�/�P�="H��;Df}�۟'��h���vߘ�Ɨ�ߓ��6@��\y}f��jW�`m� A5	I�Ӊ��+��r��h��#��:��ǳ�TY�C�j~E�����;�6��׮WxY�!�|��u]H
FL!���uS���c��$\1#2��d�t�⠀�]��W� �w�>����_�;0��6���ā����mZ{�Ŕ��vw��=��E�$7���I[;�2i��NS�9���a�(�Ԓ���� ��Bo(6�������%��iX�5�|�4V����+�N,^W}�rVdSL���wI�ڀB�q�|�W��!�N���K�1:����ݗ���Zy�V� ��E7�����d����<��O������.e��+#-}�j$g���n�ߎ\�<����߷��<%Ri��?#��OW�������z�Tk��z%'��}��s�Ջ��Eժ7W�6�ы�є�R��ʭ�th�'��f�s����\�UR�]mv��ĶT����Z����]hB$�Z�~�m�YH.)
o�0����E'�v�+Q�d�c�E��1�,���&�,�[Z�zm���e<��T8?p����D ����0��t^��%yJ��`ZV��E�*7'��Ov7�*46�����g(bi�ܖh��6�U��IY��n��{'��Ǫ�5b�����~�OI�Lr�
�!悿��j]�:�e$��&���X>#r���y�e�0�J�ۋ�|���_��;ڕ���\	�"�O���8��{�4	�9�,]���\|5�? ^���6��ӾH�H�c�:��_,!��g��S�͘cQn'ӵT�ګ{����)��n�;��m��8C���;�!�KT��#�+)�"�4{�#ڥ���:ĚE����ZQ���ua2�.�M��=~T>e��H��̂|��3���=��
�$L��N��+����\�MI�l��#��RuR�~Dڅ'5�8�𖖔<(�˞ǴvS}�����X8�{^�s:ټ��$(^�Sr4ұ�]u9L*�tI����읣_��ۙ� K�Bv�8'�DLl�?Os���d:���^%G:�R�9A��A�6�k���S�4C6eo!�m\>��ܰ������C�ڷ����_k��Y���
���+��>��j�_��O�1r\]����+�)L�P�2�*�uIa3��}�"�����\�.k{�@Ю(-}��Ċy�r�~�`|5��3��i^�SgK6��]Oc18G- �5����7/��C��4�P��+_�Ky����\�
�E��y�a�&"���U ae�H1-�n@\�*Zϧ��*���X�G�ƾn�2�����'�}b$Z�ҁ��[��+,�B<��/�L;륞
�@?�a��Ѧ���J� ����qQ12� %0�H���q�C�,[[�S;��=Ћ��d��h�/�����xd�%���|g�P:�8h!��?}��Y��:�!�ѡَX0U�'��Q�
���""�,���@�5Aɱ1!V7��D�w�P��������Iև��V.�3���c׷k<�"V�S��a��,�*$�eH&�������!��D��_�8\v�jK[B��c����7��� �h���764r�eY�џ��8΄��c�po��o�C�K2�]���ܨYvI����Mu���,��t�{m�.6�̇NىGb�J�G�/��Qz�����f���<��Ygq�- ����<���� ��$>]��?E��[�v���g�p�Ű
Q�fi�H�����U��|� 5�"�M����C�7�f��%�9|t��7 �t�+�dTYY��L�����]y�XC���Z�ݛ�����Ț�Qɲ�)�F��-����8͉�r�0}�q�K,��J�zD?~a�H���$Tb��T�r��8�gZ"�6K���a���mh(��ZV������l`���d�$;����������7�@���fxv8béSK��m��>^7݌.�>�4����{� ����j�����J1�L�yhQ'�� �2Qtr�ma��زVrΚ��P�K�wG�9rl<��S=M:�K9�'��.�nu���2��L&�Z���s���[.�3���Ȕqބ/�^+�f썘�~b�d�Be���3mD�K^��b�o[ݿ�+h1$��G0�gaC����u1��Q��T1�(W�M�Y���e�.�Nƪ"�����{�W�Y�I�����U�螭���	�*�;�҄�b�d�L�k�]{���-�!d�`u>�zun��0,���]�A���8�M?ht˸�h�@�pz��I�d�#�nv�lM��g�����P��������������	�5�;[� �#�^	�x�Pa.�P�yT����2���a�9�`�p3_b*���=̶˶��e%��aX��f�ŬJ;=J�v��%�a���A�5;^�[����2/i������7Y<ۚ����n$���U��85	����XEz�����Y�/u�j���!�=�S�{�}��T�>�n@�[UŤ8��`cR���2�����6�?��k�f�<#�0�NGn�l�>  `�-?5E��H�����ӳ3xc��Yw.z�g�I^���2:���XzY���1X}9`1&�3��q��~G7S��
�>,�j3=#�4�f��O��)���8��=2"+�iv���އ����p�o�,���(����Q�g���i:�����PD��Ѥ\!�/����"ES�>�G��e�(��{�L�]2Ym�<����
�����a�{�:ʸ�E�-���Iu��.=�����ao�wa,pp 8q@PX����ss���&e��b3���U�4��g�r�tǂW߉���b��H=nDBZ3+m�\�b7Q��S�n^M��]��#��#���܀��c6���'��ѓ����7�l]��1�$5.J�`���S:�Gp������T--t$H-�^�\4��m�Rg����[EB���|^�V���eB���e�='��NG�'62.�G��+�pns�H��K�B%�C�zT8����x�^&�1Y�TP9(�q��� M`3��d��(p�6�lz�!W���ô��"
�~�K��a��$�69��H������2�
�'�s�{���f�m�U:Z���P�o�&��\��������/jq��UC1��mnM:OHʹ޿�jʵ���,;��|�o�&�7]p�8�0Z���HA.G�c�<_g���0�x�`dX��ܝ����%#G��\Jg�$)a��!�����(V耠��C"kY�Ô.���z���E8��F�⺯\	�H9��$����愭p^0�P�?$�������گ���oX�?�Jl��H���[^���2������Q�uL�1ws��|Ɠ�*���|U�u_��$�0�v8�������W�h�j^E����]\x��p�+��'���<4�~Za������4�I(���`�v�OW�7 mE8΀IQZ5���j0#жj9�E�wz��?T�@��*e��\-o���~F�5���P�w�\�Z9?e~��\�-�2�?Yג�	f\ ���^�W��
��Y����"��5�H���2}��ťxǹ�´5����޶�;�Q��m���H�k�ln�����Nփ�\���S-Y!�	���6�=h��>4�3q�/�ް��p�ۥꃊL��y!EO:i ��/��tD|l���
��=9O!3S�i�����Jb��(�=���<a[1�%�3�@�	;��Y������ǭ�A��� 1�흕���b�mR-Xٵ4�vz�p��>�x�H3D�K3l����p��p'�4�/�a�On��ZC�y�K�\b�B��3(�eIOPJ�Q���qg��ç2ᩤ��/��|!��`��'?��������_ئ�F5]@�("¬;q����Qe�v~�����	_T�c[8����\�( ���V��'����R/T¬D��V��_`���7S�.��p�� =4In��d�6<�r&"c�w}�'��m�S�pÂ9�f��W�.�j{��p\�B�E&m:��@C]UeO��������Z��x�����q�ݰ�J��:*��JH[�����K��������HQՁ?87<�O��9L����Z��騠����^jdIg���IC�	j��D���QA��j�OS��m��;2o�j%楻
�$�ݧE��ˏ�C����@�0�"SҀ=�]�sr��IzSO@�Uɇf�+-!�ۤ�y�`�H����V<����i� ����O��R�%��/���Y*"�1Z�o@)��d[c��2<.e����SFf���J]�>yZ!}86p����@i�x�u���C�#-�>��I̗��`�Pf
M���;�l���^��k8�*�@�Ù��/"��w���<�gY�&���hy�]=�΁�h`ϭ.�F�'2��	�c���˹0J���cD�ACe��4_H�>��lV�F���Q�
���|��pi��b���t3�MJ;�Z����t����劭6�����7��W���r�H��|�a�E���/�>��C�߹����=2��eK$��	��p�p�,ٯ.��A-'h��*�ћ�2Vg�`aI'�&躒�F��XB��ZМ�=��T��!�]v3�1�C2������Ryb�����8��ES�#dnK2=X&<��p�x�n�Z��bC$�o��F ���S	Y�s�e��]��O����H����E�m}鎬��=8�/����J��/e�Bn�7�D�*��Ě@)�E�J�1Q��`(�*��#��BC�mu4�����oI*��0^�*r r��? ����a��	��ϩ�����
a�I�v�S0`�ۣ�#Ȱ�G�T��~�����B��E��-Z��ei��p{\��n88��������_F������?{"I����8][��b�@��f��h�1U�x�$��<��j'1 �ˀoT��j��%��x��O
���Og�Oa�����9~�j2D"bC�@H��KC.I��S�:$ɢo�8aE^��k��i%9��EM������ۛ�i<���#�����������߽m��g|���4�P�z�B|9%�4�(X�:^(����^���|��ip�gYT�� hT��>(��2�O
2���jU��������$Ht;Ο?�uS�'lK箸@V�U�/6=`LujA�i�5�p[��"5f~�A@y��"c��N���9%"U�3n����ĸ�+�FPWtJa�<����t^���L6+�R	��uV�������:Âj'��j�W�;���C�Q��p�`Jw�OR>wgΨ�|����,��4�Npr�Ȣ|�Yк��C�����[9L���KiC�3?��Z��qw%��Ttx�_*m�ۋ�I�Lme�ǒ����UL�w�P�9@���B��U#?�1�ZN�i�l��2�ɱ��'.԰WJ��.���0m�Tj#Fdy�e��iR��o6E��_����|G�/�t����I8Tg-�O�r����v����
�l�֜�:%xgN��U�����i@t���Ԋ7�٩K���Ɣ�41�ay��lܕg�sO߁
�����'o��6�8�b�E��H�V	����$ӄ��AکX*���w���A�m�&����w�)����!y����~���e��^0���1r�����Y��$�����%��I+zbX��B�J�� ȏ�2 ����!VG��T�L���٢���_j�cOQ'"՛�+��l�j��d�϶Kb�m���]��肹�Wx(.�~=��v��ޭ��y�L�*JHAL��u����d�v�,�$~ٴ�����*���KK��c�6
%G�>1ٴ�}&ۙ8����W�R�ꉄ����:ޢ��'I�Ĺ���1��+j���8*�ʙ-wnu������h8S�Fb�K��Z>/�_/~��68nhl�r�"Y=�H8�[�������@�՝N^��S��c
�pl<EĖA�����`Ks� f�l.��0�U�md���]$2L��94Bq;DT�%LŽ|�//5���װ�ܔ>�bfKjҙ�6p�+�EVơ���֯[O��d����I4d���N�Mτ�Y�G�J#��6���^�$�lj��+_^]���_X���G�h9������/�j"�������b	�����Yi��Z\�yLdo,h!����U*���רJ WHBibb�={/�"��94�-��Ɣ4����Y3�m,���^-���f�d)���tM���6'�&I����{Nz%�P��R")1�����w;��Ԭ��[�F���w'M�c������
�V����L���OA����Lggy�J�S?C1�|��Ǚ&���4Ʌ�y����}N�O��m+L��~}%�',M?��}�1��'Z���5�����JBz�\��RުB��;J���p��Cm]p���ϝ��9��QS��8/Q_XN���K4�g0�}�A@.��Ɋj�s��O�9n!�(G?���q�|��Yt�ф����m�G��ԁ��6aq�0��!���N!`����\y�l�co�2K���'�
�"	�������R���!�7%�rf�f���� �)�3��:l����Z�>�1�1�.[��1�-�d(���4��������~h��e��8R�N���O���Dr��|x��|�s+�Px������y�w��R��2.��@� m�|��ڜ�M���Xm�q#uo�l��w�x�k�9&Y�&ɾ��Ol,V'�C{����ώ�A�!P���/��&�%�9�d��/7fswf�KM	D@����uv� N-���F�s�M{3JS) ���f�Ұ^7<ч�~��+B:ǒ;��7��{� _�)����\	�x���3搟�c��N�t�Ô�[`��@�Ra����� F28��:�aC�u.	:����!���]��x�N�m����m�M������*^��X~h�ń7}h��Ec\�3�P}�E�L�uF(UH�Ja��ɻ�|W�#Q��y��1�n�9������ 0�}�A��9��=��F6T�A"�Sy������	���R�����x�����ǩd��9C����f(P�5���P���9558��;�*�kBݫ\��X`xFy�(mt&&�_�~b��`��y{4bp&�+RtU�j�s�;G�ʋ���Y#�K���$���ݺ6��/��"��dU� ���=��l󍴒WW$���d���d�t���6�g��w��ݜ��=8P͠b�ct�D:A��;��'���M�� �����Z\�Œbjd+4��~��RKf���	B�d��J�"Ц��4�C��hח�)�Iy�h��_�#�)Aw>�L��Ml��]����^�P'��03�*�qt�yl&��X��\���ι�xym#�Y�Q�\��4K^;��J.2��%&_-�>6%>�,y�"ի��TW��Ш+^5��hѪn���O`@+��8��a����B,����X〫\Gm�)���פ�g�������$�72���@�{ T`�}���B�{�;8���/��M��<'��9�R��'�<ֽ\�rsx̜���l@9�<|8�H[*1�x�׍i�=����bHQ����!:���J�ͨ�@�񺎯̫!�b�7����ֺ�j~̬��U�%��s.���$!�2^,Bu�StԑEnr2�B�O0O2I��<d7�W�� �I��ܜ�O>x����X��5oO��S��X='#ژ`�%N:��*](�:s�C�+��׆}�� (��ɔ�,+}�u�H�$�����y��(��(�6`��*R�o��kn���N[�z���3�~R~k����!�?I3����8q���j��+�M�;/��c�mv
���b����hLYJ��eq���^xȺ�?Y��X�:�,�$򕅢0��g� �{J/��5��4��9�鵀��}���W!���{�'��@U�
Kd~/(��
!I�]��7X����u}sps �mP�b�跛�̠Qٖ�RV����׋��Nơ_&sNl]��|v7���%]����JD[aC��x1��X���.�{�W�>��)������hl�Y����LX��Е@P�lCX���v�;�0��z����X�_�}��:yw�n�H���9���2����࠷��o���������μ(�)M�A�<�,��"�:˟�e�5j�`3���a�wk�B���>s�J�q�ƺo�ݳo�~��7��; �(�����jJm��U/���A:� �$]�G�?-�Aw�{�V|'������(%4�x��C̜�( �"R+���J#�g��L-��ٴ���λo���I�%�{�/��+w�Ðg�wVK���ӥr� ���q���p��3@dI�����%���qE@= \���J����K��b_��=R�6��F����&��8�i���j��e�&�m�Ug���X�ԛ��1��鸕~�Ka����_Ȱu�pn|�MUb嶯�γ���)})R<%X�����Vǆh̏J�z)Č�l��Ց����!0����b���&E��Ȗ�MǄ�d�](sGS�/��)!�����ߵ$�d�,�Q�v�`x��WޡBdP������]E�ͷ���?��U������q�t���^fj	^E����,jgb���x�/����'BA�a���4�Ky&��ϲ1�J�V�V��c=�vb0�;>��aD57�;�6���5���#��qeG�	�8G�ԏV�W[�����Vi�uR5x�7�_��������ɵ����b��y%�b��$��]Of�*ϭL�*�9��^���y���$���!,��� �u�\�*;b�g�c�Tr��ͥߥ(��[�]�X���0��.P��u�w�y͗9s��:�/�H1(|o�5*�!��B�I�q����r��%N�;�u����6��PPY��9�7�-��'	�s7X�<��Wh ��*'�aTa�-��:㴧&u���U���ݿ�}*)D��ۂ6�|����8l.2�r0��������)��/�_��[��v�z�@�~rt=7�2cmw�k* 2�!iON�ׯ�`|�)���#�M�Fsǲ1�H��Ē_e�y�����ug5*��nb5�Iﴸ+�ov�Q���tXžYեO���ֹT�F�-�I�l�匽������Ogľ5�i��΄E�W�~	]�i݂*Oö�Ec�\+��<��3s9�|��
).��Wh����Ѷ�.�)��O铿�L�-�UH +�[Fh,�.�GT&|�����t���qȢe?��o��Q#��d
#�2N
Qk?[���c��<+N�BNX�\�]���I ����VC��6��@�{Լ�����[�"_�=�N9'�0�����:E��&�qʮ��h�Pܑ֬�,�XP��ܲ�~k�[g3 �w?��7�!�\���|T�ϋ�xb��o<���F�������L�.�Z5K�_��'��}�M�Ӟ��Z0�z-��6���L��o��l�d�A��~/Sol����oh��i܁�QE�P�e�����U�ʲ d����wdܗ�$p���α�8�DZ��.���ތnGY�Z2+[��}������ᵁCw��hf��.ǖuZWfe6䒸yM+�)�P�y�f�n>S��7=����w�)�=�7;�)�޴�\no�O#ԡ�����e 㾸}�:���`�����J���D��YJr��r��K}ō	�&��IQ䋀��-�^�`�⿰6iͶ0{�NuI�?�J�px�����@���/�$��=���JT6��8;�;�v$/�@�SS���Stv'��5(Q�s�P�1��"��m2>i�;σ�QA)�Jϥ���Z��iH����F�:,�Ay-��_u8{�MB�Ȍ7�Ԭ��4 ����Q7 ��L�n;�Xէ�߲�mc��_6h����� /0�5��Hĝ����>!��G��s�t5��d��N�ȣ��h�f����4Q$c�]��f=�he-$�H�k�q`&��b@�P*�/ mפNq�RnF�q_8z�\���6/H�Y��x�o#[\БԨ�@�B�>�f[���J�N��n��M1%6�?���U�sȹi�������Q�X�ʛ�#�!d���8�BPc�]�=�I�:r�*{X�x^s9r����Tb��%�ޖ�Y� m
9�or�oi(� �w���߸3S��V�׮Rz�b��g��@�,���$�Y8�,c�������u����Y�n�]�b1���U�S]��퇠��G��n�#�`���g���H4��4T
L��)�nL�1v?R�&�*wP~��e�[�@x�:�2t's�$;Q�|���t���F��ACI�Q�/���L�ӟ���u&I�JD���VJC|-Y���������^MI�Õ�ƅ�V8�Ј킍9�~�C�]h����5}��c
p�j�L�Hѐ��K��I�HT#6����A���8YF̪i=�Hs���1�?s�Ib��9�8��:4܏ׁ�+�xZʑ�쥁����O-m�鏧 .����Ə3�
�i�}��_�V���\�!��X��L�u��Q�"�a2�K���i�f
	m2��E�
�pq��/�q��j��q�����B���R�i�g�㒚0[�bIف���2�Щ��swbҖV��e���唆�I~к�W�w���rZ���#��!��� 1̣C�ox�Y��K�a���P�/|\�	f���5�z���m%t�W��6����j^E�E� X^�3���Ҡ�N��E	��pxZS!��+�Vt�����t  �)�����h���u���B\ߟ�z����:��`;M�8H����g�o��{ϕ�D�ā���~���W��r��0=K&y�"���ٍ�.=+t\'d�\n<�jy!�F��F� ���C����ѵ��MH�M�*�6�٩�:2��&��	˄�[Jb�Q$Oc���A�G�3��@r?F��Z�{�Yߖ'�����Z���8�)��|3e�9ʫh�"�3)�.�5$���
w:L'A('�5����uE0{djE�k;64���@l�O�2p@G}��9*V�#[�:_W�i��rfV!!�b�-�I	��j�c�};����%�J�K�'n�����c�����K�����y�)n3閴�M5K���D���y��k%ɐH�<�6t�z5��ރ��%��*fz��J��x���.�2�Yv�<��m��$=�E�J�g�I�@2xܐy�Ld�/�b'��y!2ѩ�D(6�v%1�I��7{��U��1�L�Ђ��`̴���*s�=�u���`���0�:�A:E�a2x�hF#K=<ZY���ܛh�5��U�	�0� ϋCn-<e���3k���9wk��.�p�E��0\Ĳ㪂[��M�tpz�NYM5uu��,'R���o�O��x��R6&d��0�����@�\�����G���к;���kؔ�'ЋԎ�e9o/��>#��J�^�f�0hkf�l@�q�aR��!,��V���ڠ_~W_��v�16**�Cy=!��b}�a^ی:�Ұl+4Y������c0p��#4$�.���ޥ^٩��W��r;�}�7�G���0p�V����䱖�F�ڽ���m5��]��N!�_��n9�.0��W(E��Pp���Y���`&�z@Z8��K>�sy�JvI_�xBEI�gH�P2��]�����1��a!o�����]����jH��*q�K�F��|5à�w$�r��t� ��9�QV^r�'�;N�OF_nH��=�UO�M�IF6]Ϡ���32t�EdH@C�ۙ�鰮l��
I#{qP23�O�a;�T2?cT=�Ј���D��G~y<�݅U<=Ki;��L���BF�����|U{gp
��=�J�+1�!��r�)# 9�I�4�T��~��Rુ�\�!��##��v��-A�4��T{��M̫��DE��X�j�]G��3r+k���2�L�߆�=����?��c���@� ���w&����Xj	��?���Q�Y��\��+h5o��d��TM#������/_6�cc��%w�)b�ʥ�6�衊�j�*�{-<���Ʈ�����4B����.(��DsP]"�����XrG4��= �X��*����3�����8NLV��
���a�?ʅSP��,DJiF+cV\�n�k�ll���ū�tS��}���|�u}���b��������庙N�i��yIpP4ʰc�F	H�[p�'1�U�+���E�B�pQ�ǟib:�)�̙F�P�����	�F���P���5�ᕄ�ne)V;]չ���(1�4T�>��YyF�91�NP��)�)��*K��C�ֵ��9��/��X���~6�Xt.E\�*.f�nע��+�9@�bd��u��SՌ��U��o<k>I#�}�c4+D�_��M�p%�Wװ��y�ly;=?3!�i!ZTVQ�de��'�!zv*���壳�Z�G9%V����O�de��~;E|0P0t~e��+�kG���V�Q(F�u�]�W��KQ����5~t�Z��~Ud)=�C�3�(R��LT�Nǳ@��s���x����X���I;e�/)��%M+J���W�v3~�2tt�OL�V��d��X�"���ʗ��n��Q�{���G.Lͯ��%F��L�,��xD[	$S��}
&��Pu葭�,���.ο��_iےzX��n�-��h=H�d`��J&��]vտ�Q=�������|!�`
A*\N��@r�,�}����"سuO���_Q�t��� �&;Fm�1me��qx�nzNU\&ba�U�@|�����6<�Ro�����99[�ؗ~��#����Q��M�W>��%k�+sV*w�s{D|3Dy�_��L`(��-�c�����Q{59����K�#�|.SDf~�h�P���a�!L�yX'h\�����"�Q�^3�!7��U��t��Ϸ���U�?,�(ca����(�s�V�v�� ��:A����C��z�B�})-l��k
����������]Z7a���j���\r�I�B��0w�lĭi`&��0Pҭ�e?�	\�_��p]]���!bi���~t�s���6���@�F��T\݊�]���~�_����E��x/��Yky.���$L6�@{���nڪ
���϶��]�3~?���=_p�c��>��Q4+��h_5����wX����"4n��x݅���Ij& �w����|���8�9�a�����29t4kl��;�)_��/��T����Ou�ƩЕ~�AX\&-vt!�In6�}�Sr6�N�5���T���f)g�!���Ǎ=,U��N��v�] C��*��[��� ����V��s���������z��h(�Џ�f�"�z�$^JHKX�����!S�:�yg��j���Tf���f�4̚!І�!��ht�+�DTN��X>z�!�lqO5�v\f ���es�"4�`H�u�O���_��
��m�a�B�����8��,�����I7H9�sB��&���3�Қ=��%iЛ?�#��x�' ��Y�E2���������8%�U��8Ƿ(M�R2
��X�����`}\|���B��`��ͪ��D��)��\�]�G.��c�̝6�c���;jF�&H��h�xH�v�׺�`���rm�ח8 [ʚ^�k��5�`?����K��.���fW��3+�.׽l�S,e|P ^u6�%�܎���#ZB�y`���[�bR�Ť���� hU�՚���=S�U�S$:í���Ö�z���CΥj���>$S����I��Π4l|;c��/|�I����w�Ȩ�{�xKl)�P�:q��Y�gi��G���ߪ��$Yb���p���D;�!	(	�i�C��O=�ֹ]1C�OX\C/"p+ч�j�0�!}.��_fI��c��Z�N+���$����Y�k?�X��Ω������*p's���_f����Y}��+��}��� *�V�*�F2���K�%�&��eU���=��-g�ό����,)�ȡ�����jX��a�h�"*�_���?��&hr������Ҋ:
m����=�d�`�������0b�%0�cva��� �3%y��;/�	F�~�c7���R��,�]Vy���r��a���MJ�8(j�ѫ��'/JK{�bWRM�:o5X���V�Tde�L�Et�Sm$�2�:+!͸ᥦT�s�����I��/�A�����r��mK0���\�0vp�#�-4;;��;8�e�fcB#1��5�6:�jD��yЍ�ʩ@�P�g��$S�H�<t��f� r���y�����:�c����A����3��y�5�Վ�����Zc'��N���Ԃ�o��'�����TސJ�F~�m��f�?U��
eM}=�����Q�>\w+e��/��{�gF=JB��m3rC�ϣ�p��H�u���`�I� ��̊]�<�2��Tp'��'�a+r"���_�j#�ف��r�	�.�*>.C���. ::�}��So~%@��m��� <,7�3>��Z��9�*���!2�ΞIӯ��_`[Å�	�ԡ�T(J�N�O~�JE�����)O$�'�W*׏���X���oH��l�ɓ[T���k�^��D�F/���K\j�$�;����5P1Z$i���������\�����rٶ3$�P��œ7W�RA\���"�Le�|YU}�4��'GOZ�}̦]zz}���c�/ �
��=0��RqG����3*>@�n&j���I���:pj��]�(��]�T�_���',0����I�/ ����ǅ7Cʎ���hcܘ���(�7�&���DC��͵8b�T����)��O�E=&{��^�h,!:3D;����#�_�{��)����稬�" �֒/��ME�{f�:�n���Y(�����j㮏���
 ��
�7x��O�m���N�&���Z1ar�^��JY٠Q��R��H���V&�c�h��!+E�9r]~�� {l�{���NN\?��y5#&��W��������4E�Ŗ��Ί��`D=ۛE��4Ks�wصK������c�m����.hD�U~W�����R�n��M�ik;��{�-�3v� �%VR�Hđ�.R�3]CS��1�y c����)NR��o�P���&٪�����R�]q�D���η������:�F�Ѻ�7�5b�X������D7D�$�U�;@_&9M��N�H�&h^���1������p��s�1��$�Y�8;�fň�j'�ΟN=F�P�>T����dE}��S�N�0�[SĘ�~������7[%�c��M�m�cg�(��|IӁn%�Z*�ʙYǥV�<0m�X�\PTA��zP�&GV���E耙�A�1u��=��: �9��6�pRCc��ە�D�������g�F2wF���ڛ����<����C\�d}��ľm���tRu�,kF�	�K����
��w��tč�����{�o�����|����@\��l��d�ܤC��i0g��v��p�,��Jش�`�?��! U@7�ZNJ��H�l{5��.�uI����o ����RS5���h.�8����X���C/l��=i%��0�^�-���;��׵�Z9�N8*o������a�c�FVY��n%��e���@�ɮHMr�Y����r��<�!+�X�Y��*�16w�m�+^L�]> ^x�gd���[%��I]�,V<����t/�E׭A�WܝqP(�X����uKHLf� �7m��5��cA����K�+��-�S��&[FiM J���gp1�Ө:���c���N�8z�)�5�D���l
��	_�)N1����
@V1~~����ݗ�dR��(��E��]pЋb��n�4F�����0ס\8j�)}"�o�2�������iY��7$##��T?��X�Q7� �)��=�esW=�bwI���ie嵛�ΩIyb�������g���>o����'l��t�D�`�T�����gs��f�6$��Vu2V�;��V�� ex�ݔ�?���]%̎�������������\y���Cw/�ɻ�A�����q��d��xϦ$�q��QՐ���g��ɝҜ���\>B��D��|�X�핦qK��g�,+�h��rV���[{������e��b��:�j�fol���9Ax�{Q8Т�6m�l��B(3~ (4���/��Fs�jH�~������ɕ�"�� ���3��66���FMx+]%Mϥ �ʓWr�%#�w��%�:���Ҟ�,��x|�πLI�f�ϮOw"2��7�u�z�k�5zd�����U�>t�K���j�3[�sQm�D�L
pѧ�΋��*,t����H?$�q$|������?�&����Z+��e�p8��>f'��RTI�\s2���1v���{��������9k�S��3�d�s�O���O<P�!i}?i�4Ӆݼi��ԢT_ a�I�r����ѩ���m�m���h���Y�2y+zf�F��ѕE)��䴛V�`G����p.7�C(S���Q���mc��C6�b2��	F��ۗ
9��h�x�����)=����ʮޙY��OP�A}��`�Kz�ʛ1]W�7�!�.��<o9`	N~a�_D�?�f=�%�S�� �pg�1�6\���զ(�4�g	�`��vL�@��:�`s���A�]�v��7Med�^1'a$\�V7�]�Lƿ�+� /�5$�ҩ����9�䕙�됚����sK�bN(d���-��+t�f��{��2�@B&����A��l?�:��#���X{����(܂R��s��h�g��낆�)�9�[A8�q��6����06	��&��'#膇v'.Nk��'Y��4+�j�=�O��n4>(�G���U�`�S�O1��l�q
�Ȣ��ܛ��g�Lw>�ݾ'�$*�f��
)nZ�*E�:�(�B0��YN��a�z	p������7��	�*����j:�'�~
ܥC�	֤��/�aܱQ����@dk�M|ւQ2���ʔ�؉i��[ɨċ>�L�B\�Qg��P����r�ɰ�L+�?&L�!��b�-i�B�#t�VTh�0�#�:
SpUrI��*R[����AE��}�L��:�� |ĝSߤ3��փ[S��	�,��v�˟�-%|���ev��ǔ�6��
L��ɷ�����d�]�̝����(�/hDd��8'ch�4�`�Ir؂ʘs@v�w*پ��b!�HVg��һă�h�Ŗ;ǡj��	=���&R��Ań���Ƈ��3w] (%���Ou��޲�aqF��'c�h���8uVܮ��R��R��P8����nh��u2�A�A[�:@K}�q1nN�3���g(��=��_����㝷�����$��z�a��&C�Λ�`��I	�qq����]���r�򓊇��z�jzj���~m��z��R��u�����GO�(A�R� �����V<{mM��BaUtx)q��4����i�5�@5���s�zvn܉�T��c�	�7��9Q�@�<9kֈT�]M���v�#�ܛ�.�\i0:ɡ��f���	�Ic��u��l�Aj�Vs��`�.|�-`�%���>�?��z�7_d�J��K��is[�����A�-ga v��W��h8xw�V]d ;����lP�!��rgI=���f�̱
�"t[��Ĝ��Ҫ��6BOw�C����r|�/�o^uiy��W��AM!��pk|h#K��V��wTv���� �m�� 
O~m3a8#ׇR�G-�9bc��~1u���\�.Qb������I��u���5�^j�'u�m�>G�݊�t��A�d��LN��β#lϨo*9��'����ޞ�/�z��I��f�W�y؜1�Ń��mcz�����6i]� ��vU��(��'˴WJ�0`!l��>�SꟵo�k�rlB�����B��3�p�DJ���]QBuB���������2AX�	ϩ��K8�� i[�C�k�5�GxtJ?�6��>mI���Y ���*xi!P覶3J4�A���签	0�W����Q����3�U��4�����b����ZJ�& h�3Ǝ��J�D�~�h����D".nq����+�XCZY��k�Q����S�)wx�������Ӯ}�j�"�K�0�Z$�JӬ�j}�7x��t�B����#�(A��fD��?�n���ݹX���D,����� ���m��i��y�|K��S�3���oa��K=O3�F��&BN�a�����'�Wn;2��%[|��q4��5���)�#��AztX������g�������9 �������iA�;5�_>�����������rt��\���# !Q�� ʲˇ��=��2*+�܌f�+��z�ծ���rb;p/k^#���3T��ܒ\[E+p��^�"�ܻ�JZ98 t�0[M���%���lM�^�ʡQ�LȻ.T����L��dw��A@
WA�$p|�m��+X���I�$͜\6A霧/6�I�hE���8f��k��$��u�����s��\i�'[�7z����|ܹiHE���.	w�l.�#���.�1�T��m ��\�m��#�����
PY��[�H���GZ'�	y�W���H
%�@Nѭ�n�eѻ�a^� ���yT���8E�3�|��<"uiEրsx(��P�ы��bY�++k�X��uM�:���4��M�R�8Q�vS��!���t�c�rކ1M��Ro���_�5���pP�Gb�ND*�H"J�S����C!�<��L%��Qq��KE�<?8	!E��Z
�"{�D-������K��Y�Zɺ7�p� ��� ���&�����p`B����ws*Fb5���f��6�x<��$��5��l�G���QEtW�Q}E^����p�iB�7�\��b�O�#�u�Y���_�|�4�����)��M}�~�dw�ڜ�O���2c��`Z(&�v���30d��0����"/��ߪ� ��
���%6O��E��r6s ʺEh����I�ܯ�g��?-��T�0�؍zn�uJ��7&��)co	�Y|ڧ?<~򉘛��/\�i�"ja_�3>���:�<4�Y���m�=���hS�uõ�k"�R	��� ~ȪR˩��v�m���nG�����ַ�@��%�5T��������ՠ�h�)˂x��C�a"��#�*��6�\�G�4`U_15�c��� �J��_t���"�Bx߾�ב�z6��=)oہ���X��|��ζ�*��U7!�֜`	�aLI1������<(�"g�j�Ft�h 8��lH�+��K!�2Z�d�W���;5�S���7�*�����B�-�;Q����%M����i6�]��VX�`�D<Y[��n`�Pn&�ǀ(��*p3{��@������P�����B#��CΛRv7vS��E86�9u2��B�f��	�"
�5��ە��&mE��L�jW�b�	�{W���u57%W/�X�]�qm�G0^Bq��uE�^g�������^�Bt}�����x<�eX��*/gvG�ۢ� �[o�u���BpvB9�N�o=�\�L;��BC�}If39<#��wK�	��o)��萡��9<�W�Q���g`X>�`�X���3k`��F�N���l5�
���e}p��l���F%H:� ��83���0d9!_	����:�S����_}�ٿ���M�}�<���2RH�7�J����:��L:Fw��k�z��l�L)���2	�c�0�����'L���D$���^:�W�����ֵ�7��|Gfd@!���bۗ�uӫڢ�_o�ɋ��4w8Edt)xҞl�q�噑j��{q ��(0 �|��w�efl��Y��� ܛ�b:GGt�}�%�gV�ʦٔ6�M����!����Ә�Ʉ�\�GcZ\n�Sg&|�l�dm�Zh���Z6��\H���t��}���9�l�d&M*j�Pt�fx�k��Ɨr�AYY��V��Kare!�6ڼK��t�HB�g{Y����G��0�a�'���V���aZ����� 	g�N���n�b:@Y���t��f�*O.}�D�G@%��ݰN�`x�5���ƳP���d�C�%��y�ߋOpj�w�䠕�A�X0��B��ާ�iD�e��a�|%=v�j�ύ�>��<�#0�}V�p���Ш����u�m�}�C7��T���62��_hJlv^� 	"��uXp���C`H���O�(�9�21G����$|�j�H��a��z���)��?�u���3Ӷy�Cˠ�9�U�}�Y�w�3�&r��c|$������h��w(V-׆`���м\N����� >YDA�������
ί�N�&J�bW�4�0j�X&V%���l���U:x{��ϸ>��#�#��$�lX��D��d�O�p@/�/M���n�-6,I���=�m<���z5��v1ğ�0�.��n9������"��qλ/���h����S���j��S����@���Hs��{��n!��٦�ҿ��^s$���m�(W"3T������!#��7%Q�y�Wl�`g>�@��d�6�]�\�{��|=��+�k�:I{V�C͔�Գ��f�3׶������IEhr,��ѹ%��3��+:#u��-13�s�:^��"�SW���K{¸��� ��!"��C��)��[��!@5�uR�m��w��xPH��z,��f�.��fG8�] ����3��HM�E+���#3S	�e��s�wnv���b3I���&T2"������v�då�)8�OY>�3H?����s��
�}��Bzz�U5���Z�ׂwAS�V|1��K�.��c�o EW$=iJ���7�0�Ag؃EZ��y5��,��u���u�Ë�x�Q�E����b���e�=���Ğ+0��s�&^g��E��O��Y��Y��Ow���J��/�����z!�gR'V�hR*>Ԇ�	WBj�.e';�mS�fƇ�н��OW&�l���1@������|�!��t�h�N�@�.H̤�l��pC�M\o�D܅��X�����R�ۨ�_۠�;��Q}R��>̗?El���c��E�{C�"*~e��:&������`���ph�CAt�c��9s48J��V�l��+��/����/��8��ڣ#$2�p�+l�و��r�w��G�����ũ#4����U����T�HW��&ӈ�Θ��-�CƘ�M�<�0�P���|���Jp'j���^>�LF���&��泄���L��'�l__�BO�o�5�"����B�S�-c�5#H��:I@pNЫ�8��?R�f$ۤ��1�
��z�b��aG��f~�dY]����ϭ5�h$���� Z���:��m}�VR{��Pp��}�T��\J����
]��y�ۯ��'a$�g�zJo��	s��]���*Ԏ BI�&-K_(��_�s+�i�}��[�_��?"�!� �i��M�)0,�Ƀ���A���}jSݞ��݋�|�֑F��>�S4��HRz���k�@0�J0�U��������a۪� M��
 �H�*9�� �P�_��+|pv��LG������-J3��?y�h@LԆ|�A�8�&BN�E�/�Yx��G����K�pQ��#fR�?)��1&��%v����|�z�[�bs���`?��͋Z������|��ᡃ�ӟ ıd ����a�XK�8D���-$sT�v 6t�����S�Ե��=&�4��	���;���#�:���aCp�DV�\��=��#��yХ�n�^[<k0˓��\|�v�}� ��0�}�����Bj�i�Z�e�i��Nn=d����c8Qꯉ�(zGDJT���m�[6?ݥ�Nx'�5�,�@�`��q�$��O�&n�+��	�T��_������c�	�7�;����ݲb!r�NG��`_��k����o�A����V2J��;�%�{y䔧��o;�2�����=0@�ׇ��-X�i!�z�R��ְ�^� U�hAzf��f�isVc���?��6&�P�"���묏�p���Ng��uX��,W@�nZN��s̗�E	`'�Wy�:'pc�l��R�G
����q����>�4��+�[��Qtb�؆5֝3<�E/�¥���yz^\ˢ,�a"tT��)G�;��k[!�ݓ^�����ȳX���%;�8��e���#^�p+�
Y��E��-���((h�H\֮	ez��S8�w p�T�fĝ#DǏ��9����sB;�#�}�Iv.���b�g���'�7y������i?w��)�~Ϭ��R p���U��BB1BC% �JA�䀣��S/�vd7���[���?��ނ4��p�݈/ EA05<�S' �\$P?g���8�jgn�2%�#�	e�8�n^_o��8�@�QC#���ڢ�L�;c�K[e���"��z�kkS"PȆQ L�Yk�o�a��L'N�-x�����.#��&v�͖V+~��P��.�ut
7I��jS{V���癤_��o�װ�trbD�I��G^�BH_b"p�r�B�l��K�$~N��g�~Lu��ˈǹ����@���6�̜�"�:]�x�������Iu|�F���'\�l/
0 ���f��мuu�4���C��Q����*!z u;��z�ɽ�3I���7��� nX7�KsI�6�	��=$���Ϛ�Ю~����ײڤ;�M��ت`�qǱ���A
�1�vX�d|�3Z����<JT��qz
&�>d�|i�IМf�nǲC�=�*��zO���f�z�Va�w �+�U:����P>�8�FM�z��o�${"ۑ~y%�FtjO���-�e��`�<����o]�� 9���jV@�1lc�"1���Uڰ[Ē*�f-(��ࠕ�脎ܷ`���S�����H"�B������p�mJ�'�U�-Ҕ8����(X(���&Q�2��je���r���A�EH����M�{�Yz.�4�&��t�RX�J�M{
��#G�vPe��Qt'j�D#ٞ-�����@��G8��8�<�(���D���]�۫��k��nf��y�k�{v��&r�Y#�f�Xׅ��Oq�v�M��	s�n��g��Z�/���.
]L}bL��t�C��H���\�	�۷�au���$A�ƛ>.w�=u�]#f�Մ�3�nO.�b���*��*{_����V��Kln�Y`�	>I�����
���<- ѷ^�oM,Ȥ�YC)�w~��2�� �X�l��]$��d����Ɠ������H#Y2�Wc��e-U\D�Y�m6i�M�Ύs�Τ%���
1.Po��4�\��1�ɇ�������L��V#2!?kB�)����Y(�w�cc[;eU'���u�W:��Ve�>\����Z�=��D֐V��v	�G�J�=��k��b�w�8�an&���X� Õ���lxv���K��G N�&R�u!"w6�b�g�!ʝ����Wħ���}/b��� �]P:��0O9�b4�$t���[UQ~9R-�jm:~��ꯁgm{:��iatH�G8^�W�᫃#�A�bo8	�|#�]�����do�����,vJ5�t��e�tM�^��`E��/6�d9�	�#,?�u�`1Ţ�q4*u�X�oPlǺ��V����6d�_.������*D�Ħ����=e�(f�/�9�����F$���rq��a��}�e�%��(����]���ɰ*�R!�~�k�^�^�G�h��՘����p:Q�1�ӵ�� ���s ��`9;��T��ەZ��m�c��ުw8Ph���23,�\U�*���¢]��_�8I҉�@���F����v�(^ ��0�!���$�K�f)6���]���7Ih5�>KNIw�oR�@5�,x��]�g�~������iԵ����"��A���g�X���<��������'���s��[kN.��!�z��Բh��������#�N�	5�5u_�pWw�����ߴW*b�b<�uZ%K���j���`�V�gqV����(]K,�	 u�L����+h�#I�&�9kZ���x�dxb=���z�v�b��|*��g@���5���@����y���mV����[��Fm�:B�=ԉ��'$��C�S�ӣɛ�gn��i�Q=�j��j�Yo�x��/|zb�!��X
��j���a�88�C���p���}������E��B�՘��[%6����2�#W�7V��6�d���Mμ���+���aë]�v����[2	 p�����������n��)���-�[%zY"r66��2*����O�ƒ��]p~U��3\b���1�g�~3B��d�a��<Wu�9T���JxB.��ɰ��(�\G�����$�U�A�;ws�h�шm�-@R����Y�1���3	���y�}��c��$�ۘˀ}���&{Z1�Q�Qz�sY�Z^vOYa8(�{��c-���q��>�-4�iY4^]�g�k�Y�e�	y<����1t�u8*k������M�:��Mk�CQ��0�\��l��K��̅M��J2:Is��w=٫���Bj'���K�Y��۾{�!�HslV���qf�iM0�9sO}}���G���sj��A��m{�B;f���*��3<oƐ�̋�ւ�D��nn��w�R��Ɍ�~�>��0B3��
��$"�tў�]H]��2)�L�����g��0�!��'���£�\+4�ǚ>NC�8,��B@P���%�h5i��[�+ܮl&w3���d�;�UD���̼��Oe�$[T"�*j�W���KSy$��4eP!֎w���J�*�+t{QYE/��0"Tx����/���P��H�2�ˑ���Ww�=#`���=("���������Ǻ����au՛ ��Bxuܢ�2�3/�J�UEi�U�;��L�(��4IDc��Qj��J�f�w�9�੭�C�H����Q�����W\U�eܢ�}9�g`�F�/ǓW�L�N�ڜ4a��I�O �;�,Ƅ�9�^�kݒ d��O�g�,�KX��&5�WBt�7��(�9����&v�q`lLa �2�,���?��R�J�X�����㓒�`=�-���:���G�rI�"=�
�Ɨ�x������:_5��˸�s>��aŧO> �J���ۗϿB�u�	�K�2�ޣ��C(̉w�Ɲf$��RjwD���ҳ�މ���I�MFݩ_���U��#�%�%`�l�3�ֺzi싐�x}�'��1�v]�l�� �+`��p'&B�Z�+J�yuHv_<�%V�&p��l6��nI{h�l#.l�7�殂;�W���u%�(-����I�\���XFwz��v����Ȕ\%ǋjDDP:E�.g�#n0���3	�Ⱥ�`BJ�pђ`B���)<��X�Z{lt)���f�t3��S�Vi��*�v��+~T�un`H���J1fIKn�̨=G�|�?G�:�����3W��Ԧ�`GH�/�^%�ߵ�d읧�D�ihڤz^�w�Z�[0��1��PGi��� �e�e�sz�~��� 55�:��o�2J'Bk� 3���w�]aU���&��a�1�����~��bwv�Uf���6{zr�c�  ������g�o��'�P�u�"]��n�?�~��j�q1"�Va�xM�4���������@�+�;ЖF-��wؤ[���_sҽP�h}"*~���S
Y898�����	-#���6���h�����Q�������筜�Ɍ�ͺf��W#��g�7m ����vߢ�.s�BR�w��-v���Ude�N�$Gp�EXVL`n�O%��yW�_tE~[Y�=�YW>G�ͽz2A�����QT�hd.�( ��X���^s �.nS�]��h�s�Gۚ�p`.�$=eC�&[��V\�_~t*6��m���1��/)�1�mM�k��.��]��}Ep��'+OZOuB���[.g�!��U�yЙ�t	��3愆�-���k��k��a��MEBf?J��W�Yugp�$�!Ҿ���>��$�\�I ̤�Ү+�6:�&�(u�Y���~h��\�ψ�sd���Re2Q�Є�����|�[$&��r3pC�
�\�H_������|5���C
K��,oa���S�7��#��
dW�����d{="��!��*v�yZ��.h��-�����u��e�{�Z~�'�F�Ǖ�C�uŨ��/�JJ)	����"�o�W�Ωq���!˻�؂��n a=n!�PsL[A��x8^����i�k�����S�]K^e�d����'h��v��l�kã�3�!�۬+�VFv�f�05�f
���\����,[�F�����e��_����<'�L�Gx�V�0��l��R�D���uBʉC�2��+���:0H^s���0�68=6~��n"����T&y٪nÕ�� W��sr���޲R�# �E��I p�T�c^�t,�m!�<��9���#��B>^4�u���B�Fy�oOs>��y�)׉�i3��dGΰ�7�t�~��I���U7�9��z�=Z��;I̘�XP�ghMwMy���_}7�!;����j�hP1Qg��m����0�Xʀ���W���l0��[�}s�!�H��Ƣ�dQA�z�G[�D1�T���Q�qk��=s���h�N\±y[zI�\2����k��/��i�ޟ�G��Dk�8�KԌQ0�,g�L�����^qh1� ��!\2���-�CP��	�}��7��Fǋ=����%S�3�6߭8��i(�Z�|�������c�^��o����;9�:�J.")���&n�:)�fy��^���P�E��y�ywg+l!�p;c�|n�ԓ{)ýG{I��+�&ts�=�J�6��A�9,w�X�)s���İ���#B��"���o�J�]B*��E���_@i��Q�#��?L+6�&O���@�U�Ҵ�\K2^2 <u��pq���y� �:k��v��>�yi����'9C����<�(������qXXꡋYׂ�Z3@��>����3!m��s���W�m/v e6�c[5���Tx����R��"�m�#���hy��
��N˺�Z#�zw͘�Lr┝����A/��X��<24����>���2�ȱѤX|�U�y�߹��I��~�4;O���H'��7h�+�s{TN����hV�P����# ��ǦϬ�F�m m�;Q�ӛk|4�_�%Qwț%hSQ%u�oQ��wy�w�&ǟ�z�4*x��	m��d4��{�׿>�pˑY��r�����Kۢ��C�:o]�\�JNc�{���/^]�k���(��w�dG��~��"��gv��?;Hs�MyS�Ջc��d4�rVI|�E�$�-X*d�n)� ؟A!��܁��OouC$6Ӟ�XK�^���}�6'�m����t:i�<�r����VW	�*M����/��7i6���_I�L���C�q�����>����(���V���=�O[1 �⢷U������	�D��FyF�h�Q�P��,Jܦ�F_q<���v
�ey��o�V��LZ��R�����5/c�5~!w�[������Gq�*��4M�]�Nߋ������P��V�I W*���2�4�G.���@ޢJvČp�7$�2�P̤
7ZG~S��m�*x�%-Q���[�8�/��~H&D"�^�4U������<ˌe�T�?�����v�&�	h�^�/�{�$�ZZs��[�[�<-ir�7�����9��)r󕡻\]�.��P�b�&��,�f�=��J�"n38Rx6r1�H*"��H�[�u�vg�C8��p��ʛWo�n��5�Y�<8���V�;�q\���&U�J�8�*�����.��h'Q�f0���X#����UN��i.w�=�l�x�T*V�7w��v!��<�_ڌԓN��l��m ��{rU��.���?���Z��tےvsE�Ė�C^�͙2��,L�������c�����=�nB]~0��'�������d�uw�ؘ�C�/v��a\�z�����z�������EX[����H����?밄�%���/�@����j]iu��Y	��H��v̚����k�O9 ��hE;���{T��b��#0 @�;n���g��@�n��Я�2t�l\�x���7ڏ +�$��RUhX�E�3�hGm2�	?Sę�4�4�K�1�S>��?tD���]p�1������`c]N�5JFE�$+K��7��B�_��Wg��lf.Ϫ����`���O�EYڿ��S��z�:uF)�~���V؝qf|���>���#��p!���Q��d���@�����.7b�Q 0ݤ�.�ʯ���$ i��wz�t��� &59��(�1!�4�d�)4
�f�*�xm5)��JFd����l{˾y?yY4�æ���ؒ��y���"�l3���)]ET��v7�*�h/��C-���7Ƈ�R���n��k�/��W�sOğ�d�x*��P�"�TC�M��p$�N4��L� � #��`c׵�����ydIS�߯�3(�Q/���!��>dx�i��9۶�k� ���,D1�7��^(�Α���d����b�^�L<!f��A�MC�^¤�-�F8X�Ǿp"�y�Y�wC��"��e=���XxL��5����e�ϻ[�/Hg����'XS����zq�>m���Ce+y;�,:�� �e�"�{o7^(���d���b�����(Od���k�v,B�ϝ����r�Ѳc\H���:;��*��B�fxYǇ.���w�Y#2Z3?0�V�yΈ��72���� ;MW!,
���a7Η���{�����<]�b�v�+��Z�%(��MK�����0��_��V�*��
$�<\
H���֞+�x"���(u�I%M�ly�����[\��TH�@��TI�M���,}�n	�7�d�WBrY�2��4r��=�4��B\HN���(�s�4��A��VB����������>�.~�#���=����+���ǎ���۞�!ܥ4�<g�Ϳ��V4|�
�aX�_8�	�l��AsK9�`Ng���2 *���N�|鯩И�i��@�$۲��>3�����T����J*LZ��T9�ٱ��r�Mq�������1�$xm�X��M�@*9ΐqc� '�!�,	�db�3s2@9��G���HSB�)���+�����٦7"@���>Oz�MD�m�����W�[��:[CJLs�J���V�2���ѻ���%�p��G/zU[u���z�&l��|*��&�]��v3�����ԅ��{fہ���W=i�COk���M�+�o��^>�:2��f�z�M��n���wJ�9�2o�":�K�E��p�����_l������Q��l�C7T�K���J�W�$<X&����er'HR\��bYZ�G��Y�G����Ua/�f�����UOZ�2��1E�l��[�!��?���](t�'���ek�+�c|K#WϨ���CkEk_4����A�ö�x�pA����g2�O��i�ϛ3�"�(/1���Us8��JX�"�
"+-'���'��&�����{���`�@�o �:;H~�Ϧ��	�� �[�Y��5�9��G߃	�T��&kz߅嘢\8h@w� �g�1I*��0+S&Dn���<B��$��}��6�T��3��"x;R��R]n�a3����z5??�+S�y��
��m�&����ekBO�S�������"�X�M�E���R�vn]�?\Vl�`�G����b���Gy�Cåx�4���</=*�_�Jٸ��n��.&�0�c4G��S��l�G�t���;D�Z�U1�Hq��I�o<?��l����[��]f�t����FG��g���/�,}���2�+i���D1Z@"�q�3y�0mo�Sׅ\n����َ�H�J�6�����F�U]F�'0�Usa6�.ܖ��Q�{+Nra ���V�s2iޖ���E��GoT}�9�v�;3�l��^o�_rb*C��-������g]���;┏kK��jB����<�l���%��8Z�6%Y��/"b6U��M͘g�,�|Yu��+�K'��tIPF?�1�� ~���D�,7k�e�/@A��4��(������^p9�؆���lC ٩U�G�|�#+�l}�fT�'C�l�d����鞰���vu���ZI�[3���:ܠ�6CEQg�7	�_5���0�����ŵ�:N�)���Fޗ�G��lm_���_�w�r�Y̬ &��/��(#�@Y"@��x�S�+��f>w�o�D��M�ak'��0��/B�o#p6������'u�5a���KNF3z
//�����&ًɸ�U�'��ݓ����������rf�����bԫ]��@W�� P���Sw\���)1�@|�������ސ#$��i_M���'R#���}�kX�,�����8?Q�{���|�W�`>�:��Dv���D�f���|,&��Hy����#o�[_ '`� �E0�8�W�S��/t�nX|����+#}6rF�E��'�I@����(v�\��AC���P��\d�mS���L� eӷiO����6�K S���K
 �mYG�u��(���6�q��<>����b�����_S���~�
x9�%snͪԻ��,Ո2V)y$}|��8B%;Ć�Ո�XYO�X�\aXl+��UX�M��یl��R2��"h�a5����K��ڙ]cɹd�#u<�C�2=���\]�}�H�T���@p� � �բR�<���݄�)�["\�#�.dX̏;õ�
���w,:�q��|�+yhFv���5�hz�9��W�G1��M.���y��H΋��"�!���鐪Gr��NI?���n��Ii�=�-��� k��Ҙ�9�>�d;��π�B�?3�.4�֨ �a�,��#��pI���m?55��QI�d��IWe(�z�D>�/w�l�Ò�n<Ր�hɠg�i4q,�v�M�^�.�?Z0�6��r�G�
W����S�H���w���i��|8V8(�٬�N�R�/�|	�k���	�S�'����!S�ɶB8��J��Xˀ����ԋG /����y#3#eЗ}���z�̾X�*}'ICp����K������֩h줳��!�Y�<"�u��,�C�R���.�U��L��7���Tic���vR|7e2� Y��(H�� �X-w'&4��	ݾ-���Z���˱)���(�m��&=퍣ޜ�l�t�b3��R֥�K�D-�g=W���=U�+JUr83�!Ѹ�eԆK֡LK�nā�nB�-�'	N!)�m����uJ�8/�q[���H�*z3���(p��(62�\��/˾2(�� �ad��Dp� F� �J���Q2��yӜE��5QV��cXD���9��'�#S����_�'�8��� �ek�׃�2qz[7 5B�<k���f1����hP�~��m�K�b�B lT�*2Ż������JxJU+/w�{8X��4.�o�1��6��k����"N��XC;-[�l�!E���.�b_�xe����D`z�-�-��'��(oC�K�h��r�Y3{�`Ӏe��h"g�[?A0m�i3+0������
_�j�BA��rD�&�����d�܎��7:b���*�y���d+R�ۨ�kv�&��^��#����6�#/@���-p}�_��a�͙� ��;�E�-�c�9)N<�xA��ց�`L��v �ȟDڷy T/��&荮�*�3�e��5�<�^�������L.�W";��(��niŢw:��i��k`�gtU�Ŀ6���*�K�Ŀ�S�n�
�d�r#	�N�{�ш������}�9�2�\σ������Y~��Q���>�[���c��h��z�>����T?�%?$�${�%Agԟ��Ir�' �	���;3��*h�[�w��#ۏ!�u�ü딛O�4�Z X�"�͐��O�5H������C��%s�u[�S����@�I�1�e�����w�
~���qѻ �f(x�w��S��o/Uh��?��"|ʀNW�+ ۩N��j`aA�G���o/q9����S���.�w�j�I/㿑a�t���ɕ��b&<B���?Y	��nz����c�$D�^�����,wR��L�V���A�U�y�*C�Ϸ�������7VB�%fɄL�����H��n���~�B'��P��M������3\ -i����ߵ��$� ��9��3�^��UT��K�t/�!?�C���tKM�8�s�K�.=SN�B�,[#�yM�}�Խ��He�]��v��^D���|�Bt�4���Z��Tșq�UMVV(vb�į9��(ȻJ�����B�T^�4�0��QK�H��`^��p�����v���p���S��j#�R�ߋM��1,۞�;���E/z��13;�2�39Ӓ����R, ����^���@��Z�*n:uH�a����{�@���d�� 8�BE�^�	k������W�-�hoB��P����g�?R������ �� 윫|���g$I�.�:�u�w'�Z�Ҏ$��D}@MOķj�4�8T�f��
TD�\ ;;��Pb>�u�^,󵳛z��ُ��U�^_�	�������/�C1|":՚��h2.�f��H�PT]�ڂ{[��=O@~�P))u�3{}��1�E���w�G@3ң����W<���q��T�2�b��̐�> 4m]���������z���^ĔMC����dI#�P�?��w-�F��OK�+�pi��T~ʑ �K�Y%VI����=]bnġ����^�¼,_%Z:�+�?��]�<�No��Ҏ`;
1�";���q֥�]��t��ʺY�U'�|�؈�\���P +�j�c�;Wop���Lu�!�����u�`�pt{�U ��zO�n�.YCޒ���D_y61������dR��� �Iܗ�״$��@���o2>C7#m+�97V��/���𠮘��v�eaj����*m�A����SO��Xk?�si`��c*A#U���a�e�g�-9��ӂc[�,�OA����Q�P�&K.��\2�;Y���!�,60Ln߃��<�G���/�ڑ���!�(]p'%��ƥ�������Z���g
�h�Bxt�8`�����d1
������׎��2������� ,������1���J,v�V^vǎ4�&����p�����B��8��h^��Uذ��C�Ws؈0�<�iH�Z�����$�c@�ݚ���d~�Z�?	�#���}�cM�5q��hX��W�npmVߐJ�!���L9
�����>p�ZU�9AR��B��3�ɵt��PP��R��#�oQ�hS�Ǡ��)P��;�W"K�rݩ����O���&�fP�!	?�)�J�~��_�KX��@�9d���=�}
��i��<SY�V}��� tk�./�ٹO��\�u�"��Y'����Zւ)���
���pt�� /ɐ{��m�JM�H����8��b�l�$b�$U��i�eŤ�����PI��tAO�����e-�-rHk �I��ͨ>n����Vf���F�k�̤��Y�'su�N�����pb��d���!��G��h i4�����K�q�a��]a����|1A';�N�{�Uo�V��R[�zz�`�#�V+����l�\ĺp�$Ȳ�=�N�*�*��� 	ɘo�Y��WY96�5;������}���V�۩q�o������F�KEƹ���3�f���J�4}��D9�=(o/"p�MJ`K�r���^�����q��t�}1m�Q�zrB�2�^=~a|�pC�Թ�@�B���D�z=るL��R�g�X�Z|]�IK�MM�y�� 	=�u燆����|���+`P>��w���CL���.��Os3��N�Щ7��UoLA�*I��2�5�z��<��\~f�`%���oD�f7]Q�����YP�����˲�w�����8�O�@B�ׯL��LbȦӭEf����i85b$�G�����>�b�^j�Ql��wuO@Z�T� ^ʂvaE��P/G�GO(�?�l�q
֋Ֆ��y#�"H��Q=���������k�P�#w�����6� L��Yr�����?E�ԃ�S"O�k�%��տ��_�Q��Ĭv���J^x��z.N���)�6l8ׄ�a�*���)�����j�tN0
^PZ���ǡ[Ԡi.u�7�F�WaT�޺O���K��8A��ێ/H�@������>hjN�er�lf 	��9����Ӈ�s�1V��\h��ԗ�~ig���U^h���B�٬.k��݂��%Ci�V�㠬��{��OYBЭ�N�i�X��~Q� �q���oj�{�we��迼"�S)T�	K	�}��EA)#������t�s��܎2>aM;k�SzM�ҙ#jh�E�0+��OI�G!^�X��S���萴R�~D=���ؒ+�}���Q�Lu��.B�#�h�\�{���҄t,��Η���yVTJ���F���Ѻ�������sɄUDuxzAíNA���z�
l���sOyDf� U&e?h��"�@3����S�:c~>�B�D����Wd�h눅4T��/
��_c���z*�x�J�{�P��3�1�?uz�ǟD�=��VOX��N4E5)*�w�o�C�n5R�K�(�"YfQ�~	r�V�s�^q��\�y0���9�=��IT)�b��\9��j������d|0��;4���Y�E���2*f�~L��k~e�1X3������H� @S�׊�?�y�����7��/�Mo����H(x�f��x�,�d���"�Q�:�8K��(�tƦt◴0�UOkc�#���i���?�}7[�����ĨIE\�ͱ�c�0;a�M��Zm�=U��(��m������y����gW�I�9f�Y��
[H��S5��U\)z{�e`is�<%A��>F��^���s�	���E¹�
M��M�ٶWp����}��xY�_n�����xm�;ws���E�^3���4P�ye�	�G���F�Y�,����@��r�AmS��s3Ҽ�1��h�d��K���!�-�d��99D����"H�ڄQ�/ܨ3FT���i����B^$��
�#˺gg_ ۠Ɲ*�W�ҺL�D�]�Q��O� #7��C���5�p�@pdzݒ����#����CD���uHO��n���Ajq�ʨ�(�i������J�1�Χ�y� I�3?5�bJֽ'���jP�E�/���X�B��Ȅ4��(�iVm����w8�d�eF�6X�>�?�d٥�Y�p�0�j�7кrI�K�O�a�m��f�4��m�v{_kVNk��:(j�)�U  �C���ZC��Ob�$��Mg�!_�L	�����.U���Y3#.�hjn��9���X�b�ҙ8���n* �׿�o[���{x�[��:5:e�n�UX���XI.��	���#�waY���J� S�v��%6�=$q�&�>��NPn��+���yx��6��2^6�y��O�zR��َN
����p�%��(��]W�{�4��j� �,����U�<�6�QJ���c���e�r���{�X-%�݌򼹹���������C��?��}ɉU^��`0l�W���Fȡ�7���`��"Ǳ�~�{X�F32&�����QWq$�rQ� ߊPf.�I��r��jdϩ:Ua⯾��O��1���{f�a�����	�x'<��q~�4֙���t�K�1#k���sڔq���5���kjj��)R�
��؎P���-�����b�
�����G�J����}�ȤcW�H����D�_�9�W$���ᱩ�>��u���&B�W������4Ŵw�3�]�Di�L�0�X��=���d�p�|��G��[WF�g���N�N')�>y���n䆁Ի�$��=&z��e�mLn���D��86&J��������]�Z'Vg���} 
�H�wu�e R����9�H�&��a�PQ�{���C7{�؞_gA�"Z����ۏ����U~���t�5�1��ސ�3[5�\V���3`�x�^����r��U������"��������	��	uJ/����*�6s}'���4ߣ��Ѳ�J���h4kp���Ȳ�O��n�	���н}�Ѩ�s �<�Rn��f�\�ZK���YFN�ⰵ��������{�ܝeviI*��`'o���8D��N]MD�&��/����㫈��Ͷ�o����3���N�3����96��(,�v��g�+�"X�h3ʎ9f�B��AEp�%��;f�[Z�S$��Q����FF*B�=�V�N7e52X9���B)_:U���e,d�_�E�1��2L�ơQ��&x'�>��v�gZ�:n�r]#`��L#����K���/�=j=�5R�a.�̖��7��
hM��޴�	U�A]Y��i#��p�� �Q1A8ɩ����M"�~���!iio\X2��R���>���!��6����AO��=�jpG[��{W@�1{\��뭟כ�휩��I�&$6��9�x��� �E=��V-�/*ЄH�뛺{��} ��:��YΤ��d���S��A���Xo�g���K9�^N6s��3�˒8�����:Cj~9���\b����h1i
� tx�6�۾��xm� �����`�����m���a Pq�u�+����aY��u�V��_�Թ�eE�*�6�'�$�Y0&V33�g|���*�����,T�5��X(yȵ<��[n1PG��<)�CP�/���m݄u��w�}�^=3���{KR���Z��zx�(�V�X���x	^`�b����*@(��e���Uǫ�������5�O����^��!ޤz�TB/�m@$���z0p��Gju�zo�`Sͬ�σ���Ob�}ֽO1?�L�a��zA��	+X�6�_�A��i�b@�g��H�ٚ�͉��R�_��CU�-���������X�ܹ�7�;ǽ?*�So
��z>�}g���ݔ�0Cq@ڗe $�l�v���0I�
p"����Y�\����*���Q;�uo�9��t|o�Y�x���Nÿ庑X��2���0U(�D�X�;줢��H���XHƱ��S	�zX
�z1��hb-.Y�n���祈̰�6X)ʊ�<3N�CI� ����4 4`����ai��-j݄<��W'�5~A��$L���s�c���-1�=#K�7i`T ٮW�9W��8E�1ϛ��"���aEZ�ӃR[�q�?w>����B�s[�vxڽ�hDR���p�u���TX@�a�Ɏ"�L��wV�FW�ٲ0$厔;�S�U�;D�s���g�S �x�^�����[��=z���``��,���SPS n�)���wm�T�C�O�L� G��?}�ߦ*xKb��T�hJ�πG���2�7][d&J ���ٮ2f���[E����h2��.���-�[ݲ������$���_��B,��q��?|k[N�S��%RqK)5Y�\l"�\!��d-P�CX��c�~��Mq���~��{�!A�-�ھ����M��v]�߉��l��犗��v���>�	*�vX�S��s0��Ơ���PFB��<����
��f��O�R��L@�``Nʛ��� >l�z�,�Z��fڸM]��g���:���?!���m���`T�0��o!�d�!����,r����NχrT�����^��wv#X��q*��]B�����/���[���P�kpʹ���"����eܐ�OU�D�C@��(
��:��GLi��h�M\�DyW?6����䡍4�*x=� �|j��ӳ�&e�O�E�"MX�i��6�j��6�Н�<�zu�!kr!L�$��zÚLU�k��Vp���ߍx��
���S�HՅF;/���g�����r�d4��r���L�B.��I�)ͤ�1��B�����	o-��ܴ;��{g�Lq���!�J>yt�$�383���������� s�YRW�2��v�@A"��3�Ĥ�`�8+v�_�)@��v�W^��t�)�vn�m�IfD�K�%���HZr"/�v-�P
�pɻ�+�PL��,���*w�`{�,���yN#sijg�	��.P��ݏ���V����hN+����*�{�e���R�~F�Su����%hP5��g��4��$�Ԁ�V簬�k�\��&r�nՇ�_���k��Ty�T]�;�G����h�ڕ��	G�3{���w�R=M���2��
w.�u�-��~A���[ʌ������R��h���j}0��e��i!��N^�+OQ(�̵SR%�q�dܟň��ʚ�?;�y_�-! D���1<�t�X	�XtO�a��%�5Y��e��q�Hz�G�-���m$9��Íz�r���H�*!�tD���c�/�x��닿�	��+���-�x��p���1����Ȓ$���2��ۉl�X�Gtdב�O�E���[�1�z=��-.���q�W�dU�vU��2d��3�~�|�4�W��υr~�{_�\{~;��o��ڄ��(eѹ�qĳx��[A�e����%7���!+���� ���Y�:�����>_���m�C���\�=ױf��٣l~��q�?*?��6{�>C���6f��}�}�����{h�ٻ0�}:��m5޺�B�HB5����!��g�����f}�1����~ߵ��?�
����!-������vڱ~�i)�X���Y�c���J��FzB/Բ��8�֐-VT@�[5��i�������-�ZX���g�o>R;�-���d�f��^�-*���&'�P�`q��;7��C�M&_���ݷv'�$�����k}�f���^��B���� zw�R�r�������?�GaV@	|��g���)�'a*��q(��U�!���aɹ��BƋn1l�a�S�������̸e,�W�D��&�c;1�RǱ��޿Bgjc>��:���]3N,��p�,"�C��	�$Z�?@K�0̣20U���E��ӓ�Ym{��BeL`d7��6-ؖ���U��Bl~�è����TXis��P��(Ͷ"�k����m,"�=)�=6\���N�p�߿��r>�,y�zEEEܝl�F�� <%c�u&F�[|�-����J#�5�Z1�{fS�df�ODA�i����tBt�Ҥ�1�oNV�gkC������$!uE���������2��w���G���f�:@<�Wʦ�`�(�&�}�L�i���`������\�q�L�=�iΫOϕ�E2���+"�RM�����1�ϣ��N=��3��8/�TS�����}M�����<�$?˦�q*y3�p���Q�x��>`�)iU�[=p����W��޲M�a�v��h�1�,���r�ׄ.+�����/}F��a��${��`��sթ.�|��z���΍�	u�zbM���M4������S8����ZŠX&��D#iH
���+-z$/n!HS��&�����	3,�uE��/A���2�ٯ�F�CD�{�k��B�oi��C-�#�@oRWh�
`g�����~FP�9�A���J3����.�~L�%Mt��������rf�e�#Ï�����u��X�w6J�2���j��Gt�Ž�]�~C�z�,3�q��s�hV
2�5�=�=��!� �l��S��%��4AN���y�k���'Υ��8���Vt����<���?�-��.�Kr���^�����Y����@پfxwj�2	V��=�yV�Ԕ+yJ��M6}�.����8��H� S᪘�ף�l�6V�1xF�ʄ�I���0gu�p���E<�L�5�����W��8>tg���8i�uH�;7�`���cW"\�B���ל`x���bq���145K�_z����=r���\kD-�F7RJ��:�Snue���(���.$�)�a��ڣ�����h���3O C�pv��#\� V�i��Ht��r=ε�ҝW�b¢�S���p��VaD��<"[���l��M{~�(22��4��AYI���T./f�>1o������������5*-Om���)�$.x-�,�v�2�fRt�i~`è� %��u^F�*6j�b���j���c+gP�Bu]��!9�8Q�������I�Q�n�	)�C�K�a��*%P���OFFu(2?<Ȍ<f�NC��!W9��Z�����s�锸�l��M�����qeZa���98߫Or��l_�$��xwC&�6砷�g�?�iY�oA�I���[MGW��=NN)$w$^؆m*�;��Mt�#��kG<+	|l$wś����1ۖ�Q0-�JP���
6�r�U��n�Z�+)��s��e�i��u ���+=[�F�����ϳ�uX�ɭB���Tz{���M�����v({�1�ɬ��W�$H�j�m�O옺��O��ݛb�,x�ٖ�X4�r,�Lۃ�%,��XY�s��`��ܮ�����0c{�@��vBY{���5e?��$
�Hk/�:=�O.H�b$o[��~�&ݣ����"�/��C��\�?�����K���Ɓ�K2���� �Q���D]|����g»і:@������9_E�d�¾ci�x���F�?�@���p��_P���."���ǈ����t@Ʒi�Q��������YW�+�l1�6�1��ާ6���C[,��	d���*M]v`�>��4��H
:{l$�&_���mغ�4��� 0�����j���RY�P�Č@z��2k}��hp��^J�!�s�=�)r�p�"
�����҇�򙫞�w39g����h�ӱ��&�=/7pM-�z�˛Jǻ06����i��*��T�:2QܳYY�֩�Btb33n����쯝H�
�Z+�����x�uÞa0��a3vz����P�x閟Fs�i=�� 3��v�{(P��T�1C��L�H�����P�����ӟD���ޗ$�pM���$�?4b�6/��Ϗ�ꘕ�)��r�H~핶���ꝕ���g�| ���kld�Ö��u=�32��k�
��c��4��@>_}�"��8B�nY`�|�
'g6�QfK4��=��!�b�5����`i)\����go5�E|(�*�����#�e�:�s��Ѹd���+Ӎ�����]�z{�@����1.m��*����z��~c�G��+s�-޳ר��U������@����3%J0H�+�l��Z@;�C��OES.�ĵ����_�2�GT�����|���L(��<�a�I�����>���V����v&��86��&��&1��6�����o��U�Y]�s�ĭW^��p"�϶���$ʓc�E3�{���<=��9J���b"[ؐ��z��;\o>�4�����+)Ғ��Y���_� ���+�VyY���x�����Ө@�t�ʭ�sP��s�AC�<��	�;�# i1���j����/r�a��:�o����, Egh���rm�FP�Ui�aeTQ���\��E��R�][�W\��^����lb	��H0u��U�7ďT��ϊ����Sp���]\+6w����քzq���ۊ�{x4�7�+��������Ga���|N"���Owҟ2h�{B�.I�LAV'X����q"���s�m�iY~,�2)���^!MM�M�~�s;�]�1�f���|�������I�zQq��*��2�=��X*|w#<�g� 5T� ��*�yQ�l/�1��Ĭ���I����HPU���e��?�^׋j�j��=$�Ֆ�=+�e�U��`�N����Mv>RWZ�c~�+�M�͎���i�@k�A�M����e��	]HQ5����#�^���w�g�������KF�ԼXX�W0�t%jv�����+}�R}�Z%ک}e٨���s+}Zޖv��D��j�j!Fw��͚@9��%v�ؚ�!�R��^1��y�Ɉ�>�h�7jc��H�[�����pi��?�E��O�����p7q{ox���2�RͼoO?惤����vij�J�4����E��l��6�TD�%UȖGM�W�8�5u���/$�B'�����Se���ω���ΗDD�%X]�����l�U��1�����cw���#�1��F&�?�;0�C�N�)Y�a�/�����ѕ5k���V��4\d>I/�A/�0Z�~nX#�_�F��&�1w�VRL;�V�AS��@@5� 䋳�!Az-��f�?�p��J�`�����TK���c5��@6*���?7�iۦ���INrC��Q���BX+��Od�ih=�z�>k`�3v��:|1_��f��[/��E׎!Ǻ�~4�b}v,���P�^�y�PT�߆�4�W�����������/��	Y'61�mzaD2��E;���%d��3���������.� 0Ʉ}����*C~C�z3"�����WH�U���n��1��M��&[,e��t��B�tn�"�.�� �׸\!�����#���7SY�稼��bc5m�2�fE�nAcP��OfՏ*Jc�3��o�W6�C��g\�W�o���0jy-x��K繃�� w��N��i�+O�@��~�d�$z_��<q�-��~_��$��G�V*��.V�����!�:�I�.�6z�h&�%	3X�e���}o�+x����f��{�rt��Fh���i
F�B��@Yk@�/�Ea�l��[W�Tt�Z�s
��WQ:��gH�P���{��T=���:��zQ�5�0������gI���G�1VA2�e�]C��	���v�W��#�Ӥ��oᵂ_�*K��"��qe���ai˞;2�������MZ�\��e�wk�����ϒ�\�Zä�*�����R�&'.]���@��������'�����8�>���=f��n�t6�pF�2�t�����r4�Pg(�ݏ@�2�������R%�y�E��%���$.A<���Ww�OjF��OE�vI��O��r����5��2�A�Ao9[/�+c
ݡ�-g���]#fx�=A���e#{�S# ��q! }E+mo�=p�, �}P+�5��O1��� �!mI�����E�ѡ_�"�;`����L��@��̑������w�=S�r���e�]���诼ۍ~�c�Z��l�<�+��]H*�P�����C1�$c*��w��i�YX~d/"�7�ʄ5��F'K�'qa��b��= 2d�`B�؏�A�2ri�J�[�@�C'[;44�O�%��,���a|0��Q�ֲs�����~�H�K�7~s�&S�4�y�iC�Ղ]��O+�1@F:Gyj�̥> ΞU��5��Y{��Y>e<�F����ѹ�lj��T+�v$�#�9�F�)#�W��U^�&<���HI�!o(e�d��ڪ�5�Zΰ���h����|��#�·��oo��/{�D9q�A�N�=�N��YD�%(T� ���6q� �)8���N��B�
Xu{��E��̪�[3I��"d;<�D��+S��<����`�/��9��svi�b�RNg�$��#�z6�β�[�<
�rP����եJ�(�"�S�Q0y��K=��Z�ѱ��k��!���hf��1'~�U�%�G�}�[:��Б�0hS�;���
 _��Ǆ�E&x�.!u%�O�����Vv�XT��)OpyT��pꅱd���bcTՇ��{�N��D�t�52�Jέ����w^N�M���s��C��n�n�hC����wO���x���,6'�U��y���ʂh'�0���"����{.�7�{���N���퇴�i�l9oEO;����_��(^ &�Rn�wVM9������KP���TU�D�؏~�L����DDҲ�����ˑ��� X�5��Y��]����3Za�6��ݯZ���]�@Sa���3n/+�7��:r:�J�f�4S��(�pw ����i2#{2?Lp��t>�,���*N�KQ�ӦO�7�\֛WѠ�S'J�n;�vl/�\��#�5�?����P}�R>���V���;*�O�o+Q�O�2/�w�tE�O�`��8%������n�e��&���-<p�3����)�"���_vxB�	Z�VX�b�'w7�C� �fLU��GR>ī��\��`�
�������|��.ZK� ~l���WH*Jluo�`�����l"X����@����s�ʦ5��SA���}�+�NK��E�r�]�ѴTg���Sy��i�f/�(��q�����d'���Mw��!teY�)%��>X36`�sFZ�;����6����=��b��F�[�g�'������Q�W��\�VL8 ��րgnnG{�/�ܼ'��q�I�|#�ۄ3���p��3:3�x1p��9Q����Ur��V��;�a����K�z������$�?%��>z�}�/�f3���7�I�~/�3�2ʇ�^�� �#DD��~�oK�}v�/X �S��#�"op�'߱�搔PX,�<@��S�Y���3{A�gN����:�I��>�V�g�U*{��MݟqB�:��^��[���7�y$�^��Ƹt9�)yK"g�Y��/���^S.$QۿB!�f^#z6���,���wҚ� v>�p��/��Z[ ]YaZk�z^E�A�t�������Gi�'X�����KJa-��I�!��t�]}�Xo��B���x��Mm� 9���Y�2R�ӹb���r�J�Y�������Νͣ�str؄�PܡN�˙*�Vz�I�'�2�fk_۹��"��x3#�����u��J	��8	�>�ZC�� �`>kT(-�gr3^��ͼn�c#X����_��e"��+�U����Za�+�G_��S�js\�_��'i1@%*z��I�_�����h_�y
�n� x敼�a��QV�fNI���9�2j�.^�T���X7�Ub�nЀuk#���������7�t��2���
��{�Ǘ��7"%�?=8������!��:�\"=��]��.�D.�\�j{�iO_����^�A�}�c �+��g�c� r�J-�j*���Q_�Vr�%��"�����������F���V3{���_{�Za�-�\
�X8�54%!*~�C܀v��t�� U�6xy$WwӴ�N d>�=�����T��T����#���`}�cw2�R�پ>n(�Ѝ�ikJ-�[���Ckz��{ڋ�s�W���"�;�\� .�{�9�V<Mb�η5�����AP���i��������L�A���үG����7	M<F�S��-��P���6R72x���Y!>p!"���Bѽ����y���pLJ*�wG`#`�:�T�vk�q����SP����[%�yA�-˛���j�E�U�4�cV�� �3���|�j:�8�S��Z7��1�nNS>���J� s�~V�CVp�[d���td��#;��S�el��P�Y^���d��b���`@��1�X�����5���n��.?��~ZܩC�R����Q��4ټM��+��2�}�>P�|�(�=�w������
�E2y�'Q�8��������.�(�d���L+�����+�7L�w��H����.&����4mٞRG�N��z/��OT�ha��a�n�.4�|��hd���F���B�} QdϜ��M=u��@P�ROk}����Ś%��^	p���C�*�HR�3N?�byӧ˹ϭ	K&í��Rj�DL��3炽_ 9�-ۦr��>�~>ӣ""�cY���R^�(�u>4��*;-�Z�[<��p�{�9h�Z�+XT�����kI-=�c8<ؼ���������	q`O���)�[�@t<�o�s,��B|.�S��T"'�K��r�������bS�>��QfV���ε��CB�;:�U�߽����~��2	��A�o@/{�_Y��{��)v�'��k*RjA��h�an-���vFƾiߌ�gO[�nȕ�fs�E���؉CT�*46�8Y �|M��%���3�ɇ��@�T���^�Y�yL5�0�UnP�m1^���:ϊ��=�)ս"Ya�u�^ы0��
�jJⓈ.
�`7���0�,[��k�~p�h�T�7(ɦ��_G�<���9z��#�G�淐aԀ&O4_�����Z.�r��|i����{��ӑ#�[��{P���2�M��,8�j�ɍ�[l�R��29�d~�U���C$�� �G�������3�،K�#��/�[�&��!�X�ƩD!�����AJ���xvD�B
�	ȋ.O������"�j��T�F��0e���@_�zW�d���LbG�	6=CAӎ��#Mj"�Ԓ'������:8&��'�4y �xV�K��밐���>"q��s�y!.q�v#�ʖA1���ht�eu�%���^�H���n�v�I-�1�d�Ӑ����T�[Ƥݹ��il{������o|��[��~��� .��޾�_�V_�t�u���Y\�v������b�`����Ë5Q�����Wcp �rh�5	���ց�^{�	��=���)�7h�o:Ծg�7U�Fω�ӱ���|�@}�7�{"�S�M�Z���Dײvy(R����d��o��WL���qр�'�3�}u���ѕ�|�í�P|�ۥ8o �4�E�s��gꌇ���&�W���y��b�P&���&��F��*�]J(P������=ê�D��I�I�׆�, Og�J-_�0Fo&@i�UcP3׮��zZL��+N��4���`hϨ���e�x�,^��MP����7�~�rY���$�-0h���d?Y����?��>��b�R�"��蟴�h���
Y��p0jy�y������# ��]57�E��5*$�(�i�hJ�>�qh�*p�vϋf�G�Q��j�K�ǉ�ru�z�����W��h�_8���� ����:E�F�f��I��Fx�x��T�\u���r	vj_�,�d1}Ӑ�*�[�Z��y��l̲�JJ�;/���JS�l̃�:�OnbYr�U���Ơ��$^L��8���~Ń������L�*#k����\&>
�a��x���]�o1
��mV�;��ڎ�H�7ᒈ��Ma0婈T�R$ �����99�p�E�|4�I��R>$�_�|�}�=��913�μ��20�jL��ݳ5��ôdm5	XV�}�O" �|c���J�}���.�`:�u�^�4�f}���Ђ��y�8Z�qַ'�T1+w!����k���#fbd��/�~�x��n���\Ǎ®O���p�m��Mov�)�O���a��j���O�B6*����l$s�N��V0H�������h�
|�^r�YuQ	~�@��'��m��7Owf}%�[Xg0ʵ�&������E����4��m��f_{8%�p{��H�BBA��<��.�Q�P�Ö�o�E�T���?�U�S�ϲU
�g�n�#t!�;#`^�E��s��I{����2P����td��ӝ��K��O���uj�w"�JO5uߎ]�=v+�v�FK����E�q���Ty����<�c�Õ���ˠ@��"܏�����GY�0\�	V�fn5}�O
���5\�Q��Oȓ�e]~q]"V>�zA	ԅ��XFĎw���H��i�h�x��w_�0�GA�Z���Z�ݲ7�Ȁ����q���9S�7�O
dT�zIh!=5׿^����&���-+>P�քi�y��aU�t��;��b 	{o����1�nz3wL�]���w��TV59יmx6=�'�dF�^�5}� L�Ѵ��T�#���_c����6�M���\�gP^��8�]����B\i�ǝ��A2���ܮ�9�0����p�H,]�Ä℣�,�  �0)DqM��V�_l���ߒ'VW� _zh�\�`��낥y0�%�땘H�D<{e��P���i<&ڢ2cg���kn3-߄ �.$d
�z/Xc2aʼ��>���W{�g��� �pߓI K��ʭK�QZ>V��Ȩ���� ��hW4�Xc(`\��)#������k2F���k�B�xc��(eW��h�v�YF7��u
?A�k9�5�������M5D:t����^�f6�����^y�Q徚^Ž��\kaOՌ�ziD=]p�/Z���uDh�.�}�kz,�ΐ�i�7�/����p��iU��J�U��	�N�&�?~_����*�R�$0ͬBI�򌖭��J!1����6�E<5[�zy�<�D���:�)��o(��Z���5|��Zg	��ڕ��^�p�NP���j��EfٚJ�+�&�@��Ă�YvNXnP�ϾQ_�c�Y��d�X��P�����p�xZA�g�G<9�q�<$���[J�d*�w4��G�<�^��J�84��H�Kya�꟯*�i��S+so��@�hQT�Z��5b���r,J6|m���T{K��?ᙑG4[����C�����x<���p����S�˻����7�����D-�������k2 �8�ڀ��#��骼�/#�)��0�f �ac�����u�&�-��J�	,��8<�#��$��:'� i���ٹS���#Y^�\�sl�
�v3��TV�u�[��/`�+׋��^�nD�A�ُ�#6D��n���T�������Ē��$��X���s�<ܵ�o�l��b���M��(ю=�S��W
7z�:?��c��ql2�m�2��P]J��j�Gw���u�`9�h@�nZ�׬Ӟ�K+�'����Q9���g��z��\��|O0��O��5���7j�Ý���e!�K���)�4����VE�G�h�2"C׀ր��-�Iz�M����s5�8BĈP��T�������옊bh��������äc"�|qo���@�U�&+��v��4/$��4yN��$d :-W��dDB��צ�0��QS��I�����w��?L�Y�F�Q��Rs:ٙ���.1�n�����~���]�HC����w�3c��B�o����G� ~�s����0
;BL����cZZ[����>�1o�X:�A"fMbz��ٜ�n���Y6�z;�8(�ܳ�����wȥ)߹4hD�\¤p��2s�^����4o٤LRA���ɔ1i�)pK?@�=�i��
�^#\���}'VKo��ɭ�}���ypoq���&>-���0�Z`)���c>���i�?���4��Dp	>t"���-�9#&�I�\�|���z�֭5n��.�����i�^� �V��N�Q���Yk,���V���W��D% N��y����C��NO,�-�w�}�A���'��fO��*pb땁4����҈R?z-�m�T�������@���R������@�p�{� 0��\���Sα@��n��٭�'��}�Q���͍OGsc�ö�"*]��\�
b��q�7O᭰�����cK��� �O�a� ����}�Mil��pw��Ʒ{�p{�קM`=Y
ln�w�ɟ���אgz�Ԥ��%mb��~�J_	.i��*�|� ��8[�hE�i��%���o�k6��+�$����6V�S>A�	�n��}��à�q���"
,�:�����x�� �,L��D��֢����A�Q�U=f��|�&��(''�=�����
a72 䈺E�Z��q02�w!���i��aĿ婎��M�d�T���r~i�e��/��dS��p�0ŢF�}���I�@��2�fF�@��6 .�j�\E���NC�:�e�K�,� za� ���Ŀ`����BjA+���PZ2'��=߽�"���U�@�2��d@�[���C�,�����)����H6v�I��N�Z���eVZB�^c�-�gh%+���NNs0C�ɧ����L� �&��o��l*y7��ES��^��F9��0:�box�
+�}fO����"ʏ�PT�Q'�iڠ�,U��#��w�������DO8"�.s@��M'k	N!d�CH�,3�$�l�\u�i�0r�z��&�4.���衛u�>�� d
�Ԧ�f����h�i
��\����UUb��-;�{e��vL,{7����q�i�:%��N�R�Π���6e 3EI�}�� i��?�mo��B���P���Km5�d�yQ��B����N�A�N��5��a�IP�*�~�g��zkp�s����EC�<�hmt�-��O�Vfי��\���O���ꅗ
�ʧ�Nd$$f,�}�(^�^�a�w�|���$�06m�&��C&��2�k\!d[����}��� a{���T0��eU�9�1�聀��R�rK�����8�<pxK��j�26�7��2��!^D��&����5����8WJ�r�|~�q�g���@@b��p�m��<�}�kZjF{�
U�e}q��̠H�_I4d�>r�ĩ�_p'�O��B�,���2K���x��FQ��$æ5e��_�)��uJ��p����k7�l��Q�	�T��a�Z���[���Do�/{3��3��C������~i���6�	"Xִ��������J(r%�vc� o�aw�
�.p�J����Bh��������+�߬��IE��xc�qV��3��{�6?G�!���MR��I�"���U�� M�`"Z�+��l[�if�]5i��si�[��Q]��F8�r���OB�bi9(� x���Њ$tT��d����1>_[hj�#r��~ c�g�z�S~�85~oLV�6���3ͥ�SO�΀+�Y�(�챨�8����,i���n'��0��RW&����A���:.<��X�0�G���,ۤ2��y��*�{�Q/���Xd1�	59�p�90��B�$�۱E���+*�t����fLF9�פ>�P���4WST��N�V�u�8�1���\�'�684:��j���Fy�Y-�s1���A�\n��}U�-od$N��d��/�|g.����;�/�z�mU3�<Ч���)�J�|���\WMǁ���Z��<����Y�m�����	!����*��L�)`�C����9��&��x�� ��?�!�>���@M	B"��7qAJ ���K\�ǽR�0��ǿlY�^E~�����˚��_��p�bj ��=�u4�t�dΗ�G���B'�A��`>Q�D��hj��S�����*�-�����u���	���	-l�j�����FV�|�{��,r6��M�ް76t��.R��*��8�!Ur����o�i8:�:���wGЬ����}�K�A=��e ��UYW����E'u �|!6<&|b��Ç�iBdZ��td	�VK��U{^*�7	�D�A��s��5U]siI�\<�[��Uf7�u�yt�D"~�߱�ؾ\�8�B(�2+st?��m�GHMT��Ȑq+��U]-��c��8f8 �mᖟߑG�zZ���Nq��LHK(�����*r|&��X���L��-S��W���˞��D�u�@�G�R��	"�Dn���Jp���D���xmSf
�!L!!���Y�����Ў�rk��+o���!B3Q�Z�g�;�ՙ�fDc�
�p���}O������K��ϡG2��ܧt0*�t2��)E*WE�[ŌA�)��ɳ7^��O"7JKo ��h+�å�T{�~3��V��GZ���)�Jl�'	k�xH9Y�JC�N_����}
�`�$~�|�G�x6)���KA�K'Asmm�.KщD�Vuz{�rPHW�����9�Os��*��ƾ�w{qf��t��0����q=��󤠂��I�<pĦ"��d�?��W��J:��X����ɠ��X�0�(�M���v�P��
L�"(0�ᦰ�!@ s{�!�mP�#��]�;sc��V�#woO�4��i�h�=�_G�Hu�9�m!��+������I��1�B~��=�|U Pf�� r�n6er{'I�S�]rqRwQ��;��{e<w
De,_�f�`3e+��_����i��-]�;��c������%��b�ٕ D7��	6X�cjtz�wT�O6w����(/����pJ�4��ߛ�y�f�)m6��x��x;�]Tf�	Y�M�OM�`������9�X�#ru̧S@�[�����|�A1�$�x�Ѳ\��$\�F`l����z9{xs�r��}�{���e��ߠ�x���;���=������� zF��A�x��!��6N�ox�� Ρ�Z�OՉq������sF�K;Ҍ��7�߲���j�x����s	t�`+-s� ����"�A�縛/?��P���Q,�a�3S!1h�ޛx����uB+��y������ �ע�c� �,$����߻{j�2�����'��[ɘ9f���Sq�W�i��J^�5F+$>�j�|-g�I��;t8������gwY����mÒ�؈i��{D������2qF��$���O�>p�uB�9��4e���\�뒌m�;�L�F��e�b�X�����؁��)��Ʒ�2�u��Zھ�V�N3�#!↎Wo��F�Ғ)�Ev��T6�y磊�@r��[Z2�s��5��}a i&,-��_%��=u�⹟���Xfz�����^�>QN�4j��R�}�y
����*�{����`k��s�1�#؝|K>��̲��94xˤ.(�������ᳵ����%��	wC�(
.1g�hvF�^t.��{�WN�3<,�z�$g}�Р�K;o���O��`X��+�b�鉁�lG4^R�'4�hB<���h�"E�f0�B�v�ӷ���$�p�L��h�kw4�@d�>�"� uq��P��3��݋����	h�~O�M�˙�N�f��N�69���^�����s����i"���c `���!��& >��XX}9�zst�Ճ�
�:��l���4��0Ƽr��h��Sxx.~X�@ᕰ,�؀��=RK7P9�����U׾B�?����t�nҎ�䙙��O.�3；��ʭ9*���7��{�RYcTūʣH��(�=%�]P�w��R�_w	�C�����|��F4�R+ʽ
7�F�c���
C=1�r����hu��n�kD��,!Br��Gŭj@�@��]"���|k}�
yY�ΰ7�֡N{�eWR��>��:FEg!eI1|�&3^��77Q�b ޒ%O�����C�	�;( ���8u��ڃ�n��/'���٬F���q>R�MU�_O~�4.� �2U�-����%�e4b���:���N�5����#���4�X~������D�f��u'�P��[h�ڕf���v_C�׳��y��X�9�L�2W���b$e�9�t�2F�v�y{a��]�x7Et�����nd�ĽE�ㆨv��!�N�D_��|�^#�ķ��oa1	ܺ�H.�(�&^�bW�;1c-H�c����T�p8�P���D�W+z� R����+a3�4#�]�԰��T��$���c���6���˄��0�q�����x��T����P�D1�S�靤�g�R}����Ձ���{NT@<oSZ� 0��o�!�7����VB� -#X�U8������r��;���^l;S�+�TE�����kM	����iĺ�VX:e%���=�a�^Ew;|��j�*A+�jC�~J�Mg�k�P���P�G=�ϰ�4dd��Rΐ�d��I�mfo+�p��=+���>�.��}�I?��$����V�a�F2��"�!�����:�xuv�6�vӽ�+i`�v����ju�1# �oRS@�B�����nCsS�TYn��|�o�E��D�2O�a5�W��=��P�n���̌�����W�J·
G>
�a��x]c�ň_�o �2��8>"�a��kf�N�����֘��:O�&t?�LJ������)a��A7]^N���=�a�-���:�8��p�2S+դ��*WL�����tm>7�0�9[�q+��28A�!��h�L����G��� 
Wz��$ �z�i���=C���	��D�B@�l7~=C��O�T�5�[a\`@�#Tf�u"{~��'R�!����Q���%	d��7��Y0@��v�^��1��hb�7
(�(D�]�h��@�}CFO��n��a��	S�yT|��t9��8��'A��:��rJ_=�3z����gp����W���znO�J�� %@��4���C��,L��Gh�m���ѐ�I��;��Cmқ-I%޵����l��{<�0NR�-怸N�n ���O�'&���_�+\HpS�!ʎ6���4��)VJ�<<�r������n��q3u�(�TK��f�6�����+P�4R�q�Nd�ez*�wn��W0��~���Bmӊ���r��tU��@[#� �t:H������~:�E�i�J<��B��2�ֻ�MXC�zﮀp�a�� �%�6��+���4�f?�:��re�8"���Zk��Po��3����-R_�-ƚNn�6Ȇ,���Zs�S��T\�j�P[�$����wY�k�7�P�ڄ	f���a6����w]OU��&sWq�삖]�檿_�X�q"�2� 9���J��P���A�l>qb�(�!̉( V��]-y���aI�{��5
�|Q'��d�-�"SG�:T�PC@*4';�&�KU�vC^�-�2�k�_ݭ=�=Զ��j��&xJ���i�&��4y�ba�T��w���K*+=���c"�	e��6!awӞ$�k��Hvt=v��Q��`�E|�g��{}�zw���	c��Q�Oaw�!�W���S>L���eu���F��&3p�Q��>|���,������(�T�����F@���2��HըD��HP��]�\�P�B�Lc0��~�>m,v���#-~���xD��{�u��>�\���-�S�����nW�����j��@� �5o����L�-�M^����O�`�����S��|���(����	�$���lM8�-jA\�2n���������v�v*�j��\P�wN���Nc�Ï���D���_�m?���D?jkrY%b4�4���|~�'�I�*�ۃ@��������8�)��hE�~y0��1���O�W%>���u�����ih�y��6:;7����M6Q �h�G��E�~t�{��o��*:yf �/훒ĩ�n�(W���,�GB�I�Sb
�� (p֔B#�0��o���-����u?���#@�4�4k]O�_z��	a����%xgJ.�ۆ�}ֱj�"a󏺰]�Ћ	�:
E�njUG���wp�_D����<CeiM����o� �o.� ����7dk$趗�F9J��4ˎ�0k9��~rJY�eF���T������>ʔ��w^�.��Y���-p�����~��B�WB!��tv<���j�=ʉ1_��TY�'ќزy�'s�$��6{��4�ۀ��'L4Gp���x�����p]�pV�~�����Z�H�(�0�0�ӏ�E y ���"�X�,�b+f�߃��eGQ����F��ot*���>X�����J������?���IeO����M`6��b��M��2.��d�d�S�`7W�":��3�FJ���tF)�{8�D�Nm�Э��?g�J�7<Ά���yc>�����Ed#.m���\�!H6��[�y��d=�����$���$#��2�^!�Y�no�ӵŐ������@u���������ܡvj/WXn�Zw��,��cX8`��)ױ	�����]
�6�Ʒ.ŗ7e	��v�L&!�4 ~d�*#1�����>�Ȑ9�R��� H� ]�z�Ɨu�E��fq�)��w$L�{�65���í�����\���>��T-�������v�!����>�U��p��0޸Н�G�KR�e�E$~ʆ��ϱ 7����⨕
�k� ׆�Rd�>K�=-�³�Ǜt�ځ�����llKJ�X�O�sP���fD��8�s����4&�N!ȳA�2O˦�L�����;�,&Xjm��ͧB���+(�vM�B�4Ɂ��8T�lp���δ6H�C�f�t���A2�PB�ʾ_�F�fFTs ��T�3�\���&��,�8�c�<~g7���U�Ɠ	R��p�Zk�]7�X@��i�\�N�$�XRx,�v�q;�U�KG�_�[�& |��iOT��w$;����㜹����Ԁ*��z������ѧ��A&3h5���}��[~�h�o�(m���%���嚕�y��k���Qq��*]��Ҿ� M�S�~�'��B-Y��e��ȜU\�u��8���ط�/��%jO��1��>�pP'��^�o�b����ɐ��[E�����Q|�.ɧ\��B�__�	�9���@bl�4m*e��=�9���EJ���)�?6ڒU���>��L�4�q� �ɹ�/��/z��Z��*^�%�A�N�K%��o'�)�-�o�O˻��'�����|	�[��|�\���}k7f��T#p�z
W�1ޛ�=!�lŬJ���Kk=-5AM|�}��-����6ܮ"Kmwå$����e~9�1�
/�q	_��2�g��d�Fg�/@s�$+8u����;<��)��pF��u��oe7��]�N�hm�e'�D��2��`Yx��U@��jQߐ�+d��,�?�U^��G���񇤲?�<+ ��E�T���Ft�g�;j`߷�iM���*�ϰ ���SN����mQ��kF,����4������\�7E��������-��"��W/�:�xu��;7¼�T���8��7NJ�J�g���w�L�yn5J=f��t�j?|��m-/(��ձHm�9l��7W���B�6�1à���~B�	���ʻ�2�4mMF����d��>YGϨ�%�����#��d��&���:\c}W�΅P���	����4���y��T�-9�����J��	w�k�`���cr���S��R�fL~�|5�l�'�((�Y�v�F�_�p�k�&��>eJ�����k�9�R ��G�F����
)�*)u� ���o����ꊠ��Ѣ,�u���(`�4!2��F�Cm�6�"��9k`��ٝK�Uo׀�j��Y����YSF��cH`U����n��ͤ�3���/k�9��bUax/-l�]l��4�c}�%9��*I���<��G\f��+����:4.�d!L���̨)������:�C����sYH���:��\��-���v/t�ꋄS�y?c�ΖD��2m�ko��i�f��f��q�R�n�co�X,�-���7��.p��\&�(zrܖaِ��Y����qZ�FM2[�1�m�Å�3���%��A�?�)��i��޻ժ%+��ϐTۚ�>���'+)}⹜�mB"H�QN|'���=dA%vƞ/F�!��y؁�c�K�a$�:`{�v�r�!��J,j;��"6������9�Qz�	OC�8�#����,����߬@`� �`��%�ֹ`%U,#�5?��1�bg�=�+xVC�?2={zǓρΛ��sh�X��r	S�L���q�UuN]�1�r�1
�H�&���`�Q����X^��c�&�l���T!V�i�&c�X� �fʝBօ����0"p�V�/a���\B��ZREnqn����f�'�̑��M0�$2�h�H�QV{�`I*���Av�ux��-\�K�ޤe�\M���,gN�\�0ޱ��v?��ۣ=4�̏�|$_ZqC��.L�?J��,��9-?ve柃���Y8.��M�<i����h�C�Y��ҳ����H�,!eɤDoW4F�s�p��L�"�6x��ԭ%CR���M�sΈ������|�5#ʌR�� ,knF�F>�������c
�J��a�oQ| �x�u�]�D	�۾����]����Kʇ�̦H�'����8	�ؠv��P2e��y��qh����z�2{�ŉ�.��7O�LE�"��\��.���*)���	A>w�˫p�cY�Φ.�MZ"��I.F�D��A£ȯ�퉢�w�kk����\��#�F�8?�,'0���n6r�����k7h�.YO���&+Fb�aK��Ӳ^�;��Z̪Z
AIu�qu©�uk$��D.o��7��3F2Շ1v���=��%�E�^g�o�ȻO�y��y���p)6Z-�&Yk�%l ��<gE|��TAF'Р��̨
�:�p򹞋�I�[R��u�P��X#��G�����rE�_���A wy$��ؾ��H�ʼ��Mh3[<z�N�{��.Ԗ	�X}�/ET��qU����i>�A�U�M�y�v<��� �?�N�����Ę���jcW,� h�0W�f��GbąG 6sC�=;���}q�#���륃�D�X��e^�"f�OI��
Y�2�tH���{@ik��1����z���RҰP��)��m�v���W���?W_��i�g	��e3�	{%x�M���>��A�,+�@RΝ�*: ���DH��~{*
WO| ��ea;\��.uB��u����`\y�Ӂ�mL����i�5��X���+;����-�6AZc\��R��|?c�,!2qZc�\|����&S�Lݯ,Ab��毰9�ڐ
�6wOF�P%kQ���g]�-��|��P3�	�� �}w���:{��C��t����Sv�I"3�	~D&J<`��5�� ���`�8bs";+�+ܢ�fO�������� va<��I���� �&�ٜhh��r}J��%�!l�1 ��n���M͇�.�z|:��?f�H7���+F��ւ��6ҟ�~ͱrq�A�CH���4#���o/+O������7X|E���P�	����"�k����6w:
�<e�W}h���[싽R�M�TUz,��Έ�h�E��?|=��u��L�	��ə��_f����ǑozI�R�Fu/jr��Kӥ�d�-{:�!�x��{�gl�_S�Q����K2�	����\���L�/^@�`{H�w��q��t�Y!���4{�uB�ݕ�%\ϊ��ꐯ���:XO�
�zP�_�*�p�[6ƣrjb]�òJb�Y��W�K�����K�2�s�sN(�*���J�^:�t�"��d����DD2X�v��G��x�nCp�B;U6���w����;��{����kTn
�Z2L�+�3�5�5���3
v,��� ��h�)��ic�.It?�BJ�E��LU֏������8�������;:H1y R�㉨_`c������d�/�Os�#�1�!(q�����l���-�\zŶ��оӚ���P�@3��r-n�E�NA��5HH�jA���ޓ?/�VTx_���p��º3��h�Q.���.�m�s5�'8[�SD����œd\��D�����6=5������@�ANؕ]�D�x�$ٛ�]����f� ����H����P���<;	M��>�Y��÷�7�:��mM��LE���5���|�0�⨨��.Y����XS�s�2��R���XT���v{bgy=�� a�(5��V~(X�������퓿g�@̠���K�QkLw���=X�M6�o�U�B�[~h�Pp,w�Wfx(iy�c�L�y�M�/�AP�����K�5��)���j��2p���~�LJ�$	[��㄁"~�'�����UE䷭����J�q-m�T���!gch�g�ugq���VT��Y$���g�B!N�xe����Pb�{��b�x�M�{��� C���L6#<���wǸ��^�Xܩ�ۍ�!�lf�[b�����0��ڦؗ謌B��<�Ȋ[�d�/�2�vSe�x��:}�S{z�66a{�㒑W%��H���ޢ����nIH��e:�1�,�bs�0�nÐ�5aA��� �K�#V�_���\8A�a��;T4րy�J4��
��#K����*�����Q?�C��aR��eU}�8�Ġ���Xal��:�:>�����ۀN���&���2r0X�vv�Xa�W_��[�H�O:p��j<H�!�	�d���l]X����U�@��2G���#6��/ �H#�HϹ|Z���@1:� ��ֱ~�4M�U׿֠&������Vb>�nsA��K��Õ
0r���m%Z�� �N��S��V��i�g����q?��f*�����'�r�>���Җ�b���n���Y^�5��1P��?�o��6��Ð�aϐ�<�7�M��.�3NݣoG�B��5�PB�e"���H�����6��P�S�.��^�Ԭ�o��U!q��g��}�a�.�Z+h�td����P�4$��Ѣ+�T�q��_Ĩ�*]�0�8����	�
J�v/;�pp |�n��o/�.?z�>yH�J�a�y�F;�K����Xǌ���!��r	P'M#�D�9�]���t\$]W�r�|�
��T�U��o6:@�M��31��h4�9w<� 9�/�BzPy�e�G��6FD~�����*۰���)����k��z�e/�P��j0?'w�8��Xo�G�
�d�~͡ư��j���$g��+�U Y'����u�X�*�����y�_��G=!Ǽ��A9
�XyP�Yٞ��u?�bռ�2���u��T�_;H,#���G������?D%����|r�\`����ë^��=� ����}��O�O�E�	C�h;��r���ys&�\��kͫ����,Ln�����t��	�������lz��^a6!���`�H�Z����>*X�~�2�̃�>{��ԾKV�z�1��ѣ�)�pz`P��=�'U���ɼB�����~�.��������|�]^	J~�����Y�
�N�B*2\.T!oPcE�ttU�o<�
Q����E+���sFn-;w�L�P�S��sb(b%ѡA����>�UEROQ6�	�d���b*<����C�I`-��*�~w�	�t%�,B�U�����O8n`:}��?�y�Ǻ����8�F$.ᴢ0�OB;�%.����%2�t+1�<O� �N=S���c�j<%cC��f�4ryג��iy	��#,j�Q���f�k�7�A4s�-���s�eb/"�#[�J&���m({*���}z�|������xdf�0"���||C�x3�yZ}5�O|-�����RwZ�[37O����eEc��4�;��?~�U�!��H�U����*�J�X��If�:�W��v�{Հ'�:|����Pz/����4^ �y�kj����Y�Y�Iޫ$@f�e�i��fcxn\c;<w�t��N�-z��Q>f���i��5�Qt�tZ��S��7�R�:��2Ls�*�%I&Hzn'�~�'�����<���
j��^�ک&�0��:L�� �yWffz<NR���a�3�XP��e��{�`�*��B+�0�NŖ���C�pp���#EXkð[�'0�xՇc���\L��V��@�>#�N��<�q��}˾e���Ȧ�0���ƒc|{� ,6��L�P��
�=��o�H5� �?;��0��T�Q����A?h8�˚�>t$�h�5��z�V�#<�C!�(��]�ϴ|R�R��/�Q*�������a{@����]!����#����+)x�@��2�w;�7
ԃHqٌGo�4ea
H��!2�O�i.�R�d<�V���z��g��Z*�5����RHF3�YS�rߌ��&��(��lm��v5�?K�3���F��*��~��T� ��^F`'��Tm�@��B� u�Ǵ"�(49l�`F-J�g���D����a�j�}i/��WH���3���i����� ��6��* 2��x��m��᪣���#ΗNL��˞j��-�ߩ2	o�>y"R�c����)�A��*�$�V��ȸ�9�h��}�m�ٓ�j�8�ŗS#ƷW��_&��iZ	*��Pb�I��ot��`I�W���/���n��p��3dy����91��Ԣ�g��tv�G��(������3ao���8�}�/�gXo��LHǻ�5��׼��#�|�D��vn�ݠZv�s�1|�L�^�� 9�Z�H��<?���
�kբץ ��1W�w���кw������m4!<�����p�5wOi@#��H�SS�f� 4x6��`��=�?��)8}����mN&F�-�QT�T$�k�R����W�hv���(5�ߡ�����Cb���*�d���"+����ly��h����yx-v�/�gX!`<���\�.��#y�k%��*��+�v��K��"�	�~Q�>����I=K�'�
���7ݔm�|GR�=�e����T��Q{�aQ�`2�24���8��vm�04ĵLc{;��h�օX,�l�����7b?D���p�Q�O6�-�RA	�[z7Ad���k��d$��hf�������M���D��c??��CO{*L�b��W�y4�锧�E��d.�!�A���������3Q�9����ّM0���5��сV-�C��
�4�����C~Y޴qn�R�oV�rg= P���څջݖ�ho�e�=ؚ'H�gqh�yxh)�#	��-���\ά�bz-0����n��"	�C/����}��� 3�܊��� Z�x�Q4�s_"S�j}+��8�0�1�X�o�'/����\�]S�'@��\AR��1Y�
Em�sD�3	��W�h;�`2!ㅫ3ߥ(}Qx1�*m�L��ˡR_�*��,���Z1�4������u���>uF_Ϲ���=(Z �F�v̀�+W�2��#������0���;-�$8��J�36�\lbZ�]n�� ;>]��]���B͋[�) �|��N^���=7Z9�CVM>��u�@��L�_!��Z��uv��oS�7��W*FEz�+��O������a���\����~l�J~H��GW��腁yނ)�gx�WF��%;�m�&�aJ��L��Mf��U-��7�X�(�,�;�⥫w����׹�]�@��z��6�$r�KR�T�U��;���S�%vA�*l����\IX�^bD�±��t0�r�9��S8�������+W���5k5B�O����k�:����Xԝ�k�,��km��z�
�X[�J�2lϣ9�חU�pP�T�"D�OF�]s��l�զ���K8�2���_ �˾��][�xs��cwz��u�7�{��<�ߖ8�|��S.Q��60�no	Y}�ܡ��;!���,��l�^<�ս����'cӋ[�|^��/�[#;�oz�ѽy���e_% �/Օ���u��N���,�I��1����:� �ְ�w���lӭ�_��|<:����ω�o�����}-Dy��{'8ge���퍂;:����t���FFfe)�`��S%C��َ�I�=������ x����`tB��O��Bq�� T�$����6T�j����Q����	���X�1t�0ל@�Q��7DB0�U�y���lV��P#�A�P4�B���˦<@#[�z�
i �ST�(��n�r�J��U�+&�t����Z��F�]G�wλoh��j�����Mr�߮I0�][q�e�����&�B�~��bC~�z��xO�Mm� ��]�aT�U ��A��݀�(lc6�B�z��>��qsY�1����cq��cm�3~_��=�<W\��$�0���7��e�}�+�·��
t����l`�=�	�"'r�YKL}��I�|H��9IYV>>�}��
\q|%���5|",� D���(W_i���{�Sm�ĬЩ���6&���c��_+V� �J��ߩ��5L�D�oZm`��~��/<�`���v
[��[���އ���Y#j�~��j}알P��s}mC�g��2�y�R���_D�$v4�>����VD� �ߋ�
4��
�%���Ċ���e+M�����y�V�0g��w����}u7r�6�l�)��f���B��G�o�f��r��wX���l�E�2A��ܶ���^�7Qk�m�����}!tZ3����P4 ޕg��?����Y�z�aXf9|yT��|MW� �Pvh�����@x�2ir/aS 0v-��d�8ޗ��Gbv��-�W��i.�����&I㊕��Z�R<E/}��8����z��a��{�����l/��� �jOp,X�O����)"i��ض@+�b�$�<�j}�㑡�?R�c�h��z�Qز�e`%"��2��'�"f�IT���m���R6�nm��]�P���|m��s�HL��H�K���ZXkc;�������F�1E�!Q�f�{N"e��p��
��� 	�K/Lb���؁�T���i���SPc�bR�ĳc\�I��gWO��l�6�9��y�����{偛mK�I��H�!J7ʑ��>���?��'�h�D�"t�Qo��4�;��	X�Y��H��k{�������(
����xp�+��&����x�}�\����P}��@���#|TBz�r���5���F&M依2Uu:�-\|�2d�(�Z쓘~�U�ru�u�.r�µ;	��C��1�*T���55c�T����xɉ��/�3����&Ĺ|���,���/��o�ᄩ����#��b��kN	��ݺ�SQ�`�̈�c���߽�p����������� N̫IAL)�s�7nd�m�+��/'��|s<i�rG<��¦6��\&�;��<�J��Л�y1���ڻaDj1�^���A�瀼{�\����G*�LtZB�������,V1�\y��]�m�`�`�^3����Љ��~�Z���Ҋj=!Ӟ�� �Q�r��j�3�ߙo��3�'w������Gd�;��5��x�U7����9#/���LX"��ɺ�����,��
|[� �=�[��YS�ץ�c\�M�=�F�[��^���:�Z�'�)1n���X|o��b�v�M�
QFv�,iv��ޱ��k&EMjB�u�ɯ��m��p[�Z�0���ؾ�WM
 ����f�_��f38��N~e�z�APA����7��.}R�㒂gu��^'����h��N��HR�3X�>}印ޟMu6W�l�~�mɂ�/:b���h�g}��J벸]��r]⺉��4�"����St��6��q��RF�n:����w  �����Df�	QkRs)�;n4k��۳��t��C�rt�#~"'��3Z�DU�^r�C�H7J??7�{���b�����k<́%����~)l0�ʴ9���?2�о�B�5�E��my�<aa�m�l}UH�x��)�h��'���(����.�o�u�Y%#7���J*���������Q$�}�FVv<�_�.���DCe�UE�"R�����9
x%v��D����2� &Z�EwM����/�۷Ԁ�b�@(�{O'�|v���; �ҁKC��/i���e4�(+��f)���L�֨2���})��M�)ο���D3.k��|E.�QWID���.5��
y���p��9oߧ	�����l��`���8�:	���
H�����>(J!��%�ޓ����g�za]��{|�"o�l��*cK�7�TMpU����r���
��k/Zs(�4��!�f3��?=֯BFȣ�K�6��`�^����Z���4���6�:�HA[{�b �DJ�_�uQW�𰵘�9My/��4���:K�O�+�u`H
؈�;a̱�d%�b� ��0{���q�y�*o�c#C��э8|���u��f�P"Ԙ���ɼ_=,Q�#��6Ʌ�?y]:O"a�TJBN3�nM���{�A�w�zEs�ok>Hg�SCM������,�4�]����~��Zu������<�&!���Er����������/��$�� �b�f�͑��w52Ry�%w~$���*TU��Nm�)���	�ϓ7�bb�"lzF=.tr�����rB��⾳]ˌ(R�4�3�'��%�W�BA���������"�r|�>9 �[c����a�;`_�5?b�[��grJ�1.V[e��<�E���X�2�F�ΖC>�X�Y��������~Q�^�A�zS7���L���+2�P�NA���Yq�M19Plgp�����ܶ\�?'mh�;*\�4�HY@�	���'�5;�`A��6��<�����H�Mc}��k�m8��l�C��;/���%�Pm͍��s�M�U�l��wT��ZY&=
��1��o��� �x����)	gw���Ӆm����%P�g�}�#�Wo����zZMH�y�PLzh�ˑ�.�_K�F�\
C�.�rH7��dФ�រ�F��-n�1P`�	�XY��`}Ta�]�*u�Ä�
>�C;� �S���\��P&v�d'菶��Mh�s���E��� H��%[���Yk�3b�*�?�)mo�ɳ��$�5W`��*^��T$b�Z��vi������+��(�ejE��Vt�� }��FkI¿`���ӥ��h����~m��i����)m�iѺ��5e}�%��U�����~�^�n�xW�#��$�b����n�\xy[�{���U��]�FVD�f^(#��3�n� ��D��Y��n��[��zX;���Tɸ�����1�ƍ>��!`�鹎�W�w��Pkѕ�4)�Aӄ|V&�`A웝��\`P�;�mL�c�1�/3�
|��#�5�<���f�k��£	2��F7�de����j�DK(�����F60*j��o}u'��;���L�	�T�K޿q�)"-���O#�OD�Cc4([I>Է��M�����G�RǏ��8�Fz���Ljܫr����t��n���,��FP%����@� ����4�>�RE�q�57�H��W�����Y!4*@˛q�R�w)79�6-_�I�$��d1�_�$�mE�߷�%(�G�p����h�(�$��w�Tto,�}��A�S:[#}�;`�)�~<� }��WW/�0\I%�r��1��,�3��8��q�6�2�7���c�E	�u8L�������Y���h���-������7�m|��
d�4��Q+�ʴ-i���2��"��ͤH<��22W�����;���F'�\:`���Nqh&��~���涅��2�Br?|)Ɋ�qy"D�鴨���c=��p����6�Z�һ�����!7Ƀ�Ԇ��ѝ��@M�Qp�O/�^[��1=?�-��3�	�R4�ngg���z�rVެ���B�2T�
	gە[�#�뜇)�o����Ԡ��׻,J�kcM�o]a�����m�r���B�ӂ�5bQ���Nς�mxc�7�C�D'��5�ҕ>���}	�X�\&v%p(����^�0��]�/������
	A�8�1Չ$dL)�EO~*����e[N0�B��
�0oE��=���B�,��= �RЮ\aXy?���FJ� �߿:R`y!�k20�Ū1B�C���%���Ue�N�B����^�K����PsF����\������Y�Zi�Ã�..^���-��=���P�-�4̓�,=��f�T��Q]i�О�����-����š�7�\	�G�A�� s۳���5TQ�X�n�r��<���~H���VX �Z@4�����a;q�,��er�à��Fac�}a����+�	���X�=�K�t�2c���y0Y���bZ�x��r�X	��lx(����c0���Q*V�t@US��^u쒸�I��c�ٮPYs����=5ώ'��v//.�={e��I�����bT�1�+ޔTu����-�J��"x������A(��?����z��������,�íp� ����<��y`������$��б*^s�㱨�t���CP��=���L�畜�{������'�|��==�>C,x�9��p���آ~>��S��BEy�L�1!`��� �׳.��H��Q�(v-����(���\��,>y�X�(-�764G���^����f��ھ@�J�Mc��id-Uߖ����l(��< h�#�fIUC^�wB���dZn�9�.����wu���I~_o,A&^]��A5���v�r��|D��F)�-jxֿi/����ȝhɅ�F�_}���m���5��S��O��g�i˞�9�+�K��zV#���)�r<ǚo_?�zZ�Š۟�N� ߪ2Y�(f�ϕyk���M���`�J�5�U1�ʊ��|z2h����z^�������	�CzH��{r3f;�\�5�Z,Q�`��ZWz-due�A�SA7|�-`���R^QZ�r󡞽���H��a�<$A� z��k�� �! ��.ٚ�f�U$��̥ɂ�^���!�N�� }@�3^m��!������u@�B�!�O=���SG^%e���Cy`U�&7[��C���˖�wb�zP�ʊ0_�u� ���,
Ǘyg�q{�&}bc�4&OL#՞�m� �L5Ch)�	��G	dc%���vݎ��l�R�K%;��f^��y1�`��X�5�@���P�A�>���@؞�(:�CaŀP�lH����6��{FA�:X��8Y|7u�ln<Eiqq	n����/�,rm.��7��)���VQ%q)B��v6�b�P��s/�\�)�([M�� p)�9�=���ٱg�ڔ��҂������O7�;G��ڍ�7���՗<�)��~V�1Cha1�f����&1(yuN����.�����4;�Z�>]D� �,λ��h �hL�P�P�3��&p�!v��{B����E����з���\���CV2k&_rc��[�p�?��*�QU��T�W���؛�Z H��T�%�����}_{т-҉M�[�,�x�~2�p�5�:S���P��Y�&}����ɶ����[B�����V\:}�q����Jn�?�� �d
�5�$Ud�'��LW��=�$�9�)n;�O�u��)�R�����.�p.�I p�?��`��QJ�÷;�di��pٶ�l�d�B�)�I��ٍ�06A�H�Gm'�`�|��@����i,����+���� �S�J�@��JV����O�� ��
�?��o@K]_�]=��܋[�
j8Z߫E��qD��)@�T��x�����.���� >R��?m"��2=,H5��ϗ���SLE��0�%��ʢ�7���U$��6(��uJ�����q��sa�����3��:b#�<0����k�V��i���Z�?�
��ä�)z)��?X���&CoD����g���Qj��n#rǺoA�I���p�.~Zؗ�X�菞�灈DZfQ��%�ʾEq�@�<�z�M��˹�'26͞\vV�t�*6��P!��aT�X�4U#{=����#5�l f��@�b��҂N�[��ʩ��x@{wx��+� L�1���%V�`��N^M��߲�
�@�\�bn�x�Sq1�%ٌ�,g���[��}������fO�3k��S�>iϤߗki���\����D��5��;�8�%[��%-�$)�g����	�����Ƙ�Ot'�IǠ}|���ث�͕��?��������#�.�;l�s3�X/D�Q#���_B�Q�7^����7IvQ��1�A�����	 fc-�ǟl�4�	�?�1����f o �ޥ���M;?�K�\�󣟈�=m7*��`�9zoi��15����N_����4�����(��g1WG�i�_�J��YQ��yAQ�d�6=|�j y�ɖi�-+1�\�32(�h���j<+�Fw<i�9�k�@}�T�.Sd�1�x_OY6�B.�;��MK?=`�/<� _O���]�S!���ps �5��s�"�gP�~��-������7��F�0%6~ ��O�F_X3��Њb�
��	?�h��ox�" ������8JHd4�5c햫���2��O�䶷BVW;3�������ຳ����,De����N�&�Q���]���3�2W"¸�x���\�$��c�
10�i勳E��q��6�HJ/���Кc��v��F4�Ci�����|@7g�u����EC�h�<�ce�N�V��n���Rz-=��L�L�I���R^���_�{����r�����4�q�@��?�BsB�G�/��u}�;r�4�'��K�oEY6����ӚWn�l,��\�"�~µ+4Y�!�g�U�`{����NIV�L�}�~����~�l��Ed(1��)�<��Q��eH�<[4�#-���}��{�C��Vb��
�$^\U{��z!�R�n�aa��>���`��V��lٺJ#�����9�����?pn��c���%��պӷ5���#y��̟�aO~�+ǡ�)���f�"I��f��_�A�l��".�}���ce�����WE%���"�7��̰EhR����v��paL��?𷁋1*�NѦnC�ݹ������`���N�q�M�Cs{<�nK!���H�}w�;�����?iI�Z�*JJkT��L��f�VG���aY�8(;���l�[�]����ey�%(d������>�R.0y��o�d�ә�C�z���e+"R��߄�^��u<����~���9oTD�D
�>�p4�e�4�F=����@�s#�(��a�u���� �!]�+|�3E���w�R�^�qABE�o��(@���yA��������	�ɾX���$d}�\��'l�U����6D	`���~��~g>\娇p�������)���ZS�QtȰ��[�+��7Ap$�������$-lNN=��+n����ٌ�~�;�sn��ߚ�Y2""�i�^(��F$a�L!$�
�B�;~��q.L2�q�2�j�X�j�ko��Z�����X����E��u�ݙ1�?b�y���Y��1je��)��؇0[A�l��Ѻ��}��'xQh�^��roa@�͢Y��ZB!x�b�)�[S�P�*aG����4]�~3��X���f^��#��/���x}8�&*f߈���e�
t�6i�+Ξ�i�7Ī
��#uXJC��u����PD|޳����dČ��_0��⇻�
Tܲ#��]��p(
�l�EE�u�K���yz���i>h��I�2̗��\H�
���OGz�1�¿���I��TDN�U���翕�Amv�V&�D���ѩ����Z���pT5�B�r��V�����8y�,�Wr�,�G���u2=����5��}���Z,ҙ��Ҕը�ͻP���u�T��Ԅ�v��z�̮|Ɋ�lH.���1��P_���1�	|���m����r)�7>�/���g���L(�u�J;Y�VLH�u��~�I``��ʢ�6~�w~L��/����Wx�tZ�����ie
8�Kk�!�r[i�N���v��k��#c��h9Y>��\1��՘�Bʭ�ڸi���5��I���-be�z$��A@��ֶ���������ʟ��<���t�
Ȣ�!�i�^2�@G�}Uy(Z�v ㋲;Ou8�K������~R�7%���V�[7F0W.Z��,\��h��E�ʘ��6x�p��cL���1}	c{	�jH�Պ*����g�����������2���e�m
���9e��m��e[��Yk�Crv�=W��>"�	=�G �����"-RGC��C��6{&!L�B�ڼ� �����z�p��۬C��{�T��oz>�1�-��*s��X�m��^+����k�
��j����52̈́����/�*N�'%o�N(����ג�E]��K�`�K��G�h}��w�Ȼr�@����7���כ�y���/a���LCj�5�rFK�O�ȯ��5g[gZ��p���jf<�fPf�EU�H����L�S������ٟ!�z�ͷk'�c2ΒD��'�X�#��/�F��ն�u�)�ݖ�݀��E
,{H�X �%��Y*j�j������u��ќ|[���T�\d�h�o��o1����m0]�Qm��p��Df���cuaBIb� '�E0 �:k?��'��P�$����gT@��Q� 	���^pz�ڥG��nآ_�-
"gVxb߈�SL�ͳ��h�6��WȀp��Ѽ�aն��)��D�%���g�%�KƵKX
:��?Ir��	j��?'Ό;�x�o���Tȟ�4��߸7�S�@��W�O�w@"ː��*`��FD��HΓ~�4,��6����3����?_ �*���W��d�pzMĮ�0����8q0q��u����y/��TВS���b

g�Dh�j��jf2`V�h�9n�F�։�t��o�}u����n*ѐ� o=L���y!#�b����s�@���;6�Y�Z�I!�;��E�N=ٞC���rX�ZGM��pg&/�3��2d�D��ؘ%o�2��[X�*�]E�-�j��<M�Sr[�>��{����0�J����b![��	����%���#�d���@OR-���?ǎB�J��zk�qvP5'��&J�à�d�Ǟ�b�kw��o����+������\��a$�,���:�`%0Pf�v�1?�Yы՛�U��!�R��V'N�m��[w5<��*�{y�}d����>�pјD�A�GA3�?�h�Y���Ve�!�AY�v����� I��vT}ޜJ6~!�����"�ZP����P�eJW����m�)]�G�b�"	�����Wy��^_��b�{�,���:�A� 	��ە���u�YG��/�@`�M�~H� �
�Ť�5q��Ӟ�pHR�c�#����z�Y%�i��,GX��m˂�GVo�}&���@�\��"�@�3sDY�s8��Q���h�S�kS�{a�+o�x��`�mv��EO.ų?p2w�dՒ�N�|i�ڰ�>�FkY�y����%�$��u�҃��l9���*N���]x�dq~���O{�����D�de鹹`R��O1ᨬ�����r�|ve����>���R������/��0:j�!�}��'�q�����n�r9i�H>�jP�ƘRnZ�ۛp��]@S�N{��RU���z�rp��Ӯ�U�ٶ�-{y�2@�)�:�7��.Ͷ�ReH���0J&�ĄF����rM8M����n��v����ڜG �f�t!�Қ�L�"��-�����N�m�A%�ᰖ�"�*-���ó(�c��# ��±}yܵl`�&�|����������\t K�۵��)^m�kqb� �L��?�Sp,{G��g�H
D��;��k�vr�Ld5i����q�Ye�y	w|5_M���b�5�D=�ou�D<=�����U���|7�F�z�B�/����:����b�Y#��t嗓?�[Ô���s����k�C�]��]Zy�e)?�Aj4e;��:���{)Ԡ��]��L~�#�i'�e�b��1p~�Y<�qJ����MŬ��A�=�̍ �EzC�Q�x�R�����o�WK�d,����4��b�����g���ůM=ݚٸ�	&]hx`�C]Ԯ:��������D�_y1�YFN�����CH^+�)Z�� ~>�>����^�o��9��&����Z;H�yPD%�)6j������-�!�e%�	et'������[� 'sA���x�I�eI�~-L������E���J��.����Q�<f����b���(�IA�K!t��R���������B�T��w��@�*4��j�bl?h�����{�V�+�ִ=A��4Q��N`���}��=��Gs"R�ߥ��W:���6��+��񲐬���Fp�xQ��v�/�����5tRX,\�] �b]ʨ#7�H�g�m�����z��u�"��5�k.-J'%���s�j����0���:S����e�+T��7�U �fm,Q�t���D�q�o�M��J-\�GG�KCx��[�{g,�}=A��nZwd�Ȯ��eQm=�k���ɳ5U�%��.ѷ�G��2��0[7P�E��-��T;�2����Cfa򺑦+_��)V1L��G��S��9��[�CY�J�1�������ڳ��E�5~� k��6����3�'Ɖ���י0��L��92�v���N�.h`���]�!g�G%�4L�t��A��F�r~�V�X?�"����oBL��`w����>\�ي��^+�:��GT�]�����iB�|1�7����,x��{��K7ɲ��q;?,#�a�[�U�R��냍����W���N�8讕���Vg^�Ȁ�IH1
*g��5���x��S׌�h�ٗ\�*��&7����S��f����κS���������|��qcd0�G��4[��ꞑ��R�Sw]`)Xa)Q�
@�� -�c�=u�o�G��D��� 8��Ҕˑ�s.��LD̓t~a�)�ޔ�qN��+uU�`j��e�s!F����2O�UKq���J�xa�a>s/,'CԻx,W{�������K}5	���v�A"� ���+���' �H�I-�"3���&��S�N ���M	�Pn�ŷ5�`�|x�d�gu5# )�Y9��I���C"Ţ�d�����Mm�9�4��P����zg�(��9N��O�Ւe͓?\C�P}?�n�Oo�Y}�p�S)Om>! �rǰ�K�}.��\�ږ�SJd�_ 'G8��E��ȵ�H�H �	G�@���nfh�̪ݰ�uX��o\�e���(�p?��Z��S���G�����7[Q���/�¤���>0�4<�xR�W�f�`4Ry&��#U�J�Vs���He�QC���{9�mr8�E��ҫH ^ă���8�K<w#�e��>Go͸/�=�@�NBGJ=�^�:�W��[}[���T#��Ə�W��j1�)���y�D��b��6߷��iz=�$���Ъ�vJ�_��g�Ǐ)�P������1Ң5/}`��\���R��O��'.<�L�!zV�î�^6J�ѣ�^᭶qm���_׶�v�ʺ�]����K��(-9�J�"(����(V���t�e��BD�"$�p
x�پ0^��"V��&6Ӽ`;&�������F��0م����ۈAx�=�ɟA�#���r���4�M��:�:���^��P�	lXr=WōI)���E�Nk�������'p�Z��QI�%�k+2�W,Yս�-���oMc!�:y9?*b=8[�D������s�F:��#z*|E����ˋz}���\�	���ҌkA��ԣ|�4��g [pwY�m��?����}f�J~�����l�t4a�,���}���^x����7����M����#���N!�Na�~uC7���>!b��C��ؖ���IŦW����i�E����pم���;̗$Y,%t�]���/�,��$�ވcvp�nG�_�]�*�vȌ ����'p$>���H���Aw�P�O�M�k���W �迗n�Wv�'�lr.�վ�}&�_'��E�Mo���n3��`q?�lYlZ1���k�<4��i�����5BG>���?m`�f�{ʨjw�a4�O�Z�L��,�D�*-��@��5�� zz͹�<��☙��3{�l����Ԋ��0F`�{�p)#&�S�{�d����)�3<޼��r7�\ zϓp��PE�����ۄ�1	��$�⻐�'�m�U�s�+�a��y�tw�^�<c_�u_
�����3��*(�scg|oZ"MD�������w3�跦Hr	*�}�/Y��[=���I�?���:o���nۂ�7P4���L�p�z�.r�,��͋I�9�H_q�A����>g3�=����vو3������6u����2�(o���<�l�v��]v��˙A�*[Ƚ���l�EI?��O�Z�h��.ʽmݐJ�\R���3��[A���7w�]�)ƶ��8
h�!�ϠӐ^� ��~���/>��89z��� �Ao��j���7'����n_=E{��q(b<˴���GA�e�FU�O��M�%�2u�����Ʋ���w��X�I�񥑈�)���8цQ0����~ta`�.L�6)���2;�$t�Y(��[G��VƐ�'�Kz6<H���h�oC-i/�Ud7��Wj�M��j���Ћ�a؈�侙�ӥ��x!��IIO��h{T�m�3Ml���6��h������GS]	.�l�����˜O�?$�i���C[Uo�+�]QqU�h|4��^4��=��m9���j"����`�f)�n��p�}����ט�Ϸ��c1���"y�[��8��ec��;#�Ĥ��v���Ê�m�d�Gr�i0����l]�eЮ�r�r�2��X�;���F���ϼ����$�$۸����^4�U�	 ͟���Z�s��q=�6��mQDR��)�SҴ��ФI�u���ב���=s噳m�xS�4��fJ�!�S��0�{������&��a�wǥ�*����Re�8�G9�~�)�K��3D�I`�հɂ�
*@�P���6�زxk���{>�2C &*ܷ�}��&K&��z��0�V���o��,#�B6��uʮesq(�.Zw�S�F��c�|�دd�Cl�o�!��P�v77�A��L�Cx�Қ@Y=�`��DIz�
��;����;�5[1`�]&�k�q�^j//��{'|v�#��/�?��m��#5h��.��~�{	.|3�x�gO7��7f�)j�|�~��v�����oR�������8eT�D�l<L8Y���ea5�	��?�a���¥K�A���&R��ښs✅% �`�7�]��m�-�9�,�yY�?�Q��᳉P+]W��@i�ҟ_5bg^�L=��V��}̣��2iC����"z_SS������S�U�v��r,%�s�$�1!I�1	���>`�W���쉼\�X[.2��(9�eԴD�8Yމ��y?���P$�0A�s�1�~���޾�	~ga��H"ϭ���P�85����+f���F�o��o�����I�3�A����i��%�
�p�T-��R�-���M�[-y�E��N�v ��o���*�B�׺��JI�fs�J~�	�L�9���5�L��c��@�9b�t���;������ 	M)ۍ���'"��z�J3����خ���
.��aRc��h�8�K]/Z�+O���V "@_�N�@¶�w���Z��I��� #�G��=p�p
���W�����nha+�l�d���c� ���H�Q=-�N�7�iS=���&��o7��e<����z<�j�D*�D����i�u(\)*/�eť�'2��Ah�[�ֆ��L�9~\��+E2��d\{��lt�#���+�Q&�423���n��Ҏ��:���}}*�q���6���!&��X���6h�[x6��Y�%�4W�q"�f��S��q��e5��m����Y���h�*��������|�v����k�W�,�+%���=�J�U���+^�؝v:#"<g���*���'.���+�i�Ty�H���Ӆ���Z4sP���GX�0�.p��od�^�#�R�8��]� r�����<����;�+ԉ,�
㺀z���9��9�LM�`�/<ƍ�?%&!�3�`� ������^*Ҧ�BD�S�u�cǈu�
P�o���vx�^� MG�}�Nޡ�wR2n�-1������W��)>��3����d�e����@F&�/��T"�z\�/FښN��K�_9W����C������ꯜ-�r���@cN�ޭw8��߶�4rrQ��b��~����h�S�eM��x,��hT��Z�H�k���y����&��F�Jw��$mp�MxUS�v[(�떥�7�c��N�,�۫C��DZ��4��������t�~�P}� ���ߺt��{fΞ��dB��b)٘x�߶	`�PH�}@T(^���p��qe)h���8G�t��RF���Ѷ�/XC���š]�;����k�\�m�R�T�����W�{���^�ET��l������U��*��b������ȷX]���u��QG�7�*��֕�w��\�;?j�����*��� �jI��\"�X����#�_>�JB  (�DC�d1Est2�����]�9�U����3�����g"�p���+����^#�rl�U)F+I�*�Z.F�v��($�j�:���@F�N���
Y�_Ǹ`@��0q��̡'�O�_�1��"�
��?�MO�U>�����,V����P��յ�;w}��N��r�}z�X�ڶ��`�TC�ʭ�q+?WR"�q��]���V��sZ�u4Hxii��mZ��֘_k�d���e��c��ڂe���94���s���#��S��-�/wo�$�E�����a�D
�Rz<O����<�{�g�x&ޠq][=)�:YB(WU���!�#ԆOMI��ȅ}�f�:��hsr?�zrIe��tA�	���!X~I��]HqA���5�6t��os;nD��Y����6~ך�d�ݜ8��6�Q���/��-J%nFh�fI�Rs������K��|^��LE �������c>$ $��/N�%���Q���z���V�pc=@�M&��ͬ�ۏ�_��!�N�}�!So_)+�<�7��r)�iyE��L���P�R�YH�L�*gy-d貄h�O�\e{g�{��V$'^�z�F]�D�|=�j�A(�+������qY(w'C$�g?�Ai�1"��3�"q�t��X��钱��ԯw���X�z�����ۏn�4���{i5�R74�Ѵ����ɟ燘n�T���"\T僔��{���C���].��;/��d,�pD7� 
�UGb�K��1x� T���x����B9��q#�!z�����s�����⹔g��C��%�`Y��o�]�I�����J��Go
M�A�;"�#ƅ�3��b���	�=�4b
ɥ/��U�Zy�z��Oϧ�s�*!^�Rר#e���$�=� �jȑ�ͨ�93(�<m�0�Nv��FKv�؎\��K)%n�����V�R��;7���?dm�`vi��ѭu/�	�,��{X>N�Cm˫	�@�<[��z��\d
v;�����ӿ��9�lQhq�Ev� ߢ�9��Bʎf R@FZx�k�H�\q�zÆM۹NCjcWu��cg �yxU��3�̧��3���V��������W,�����+��}�d��
�Od�%﨏{D����lM�fʬ"��\��������Z��0�[���B��/�t���F����-r!Xs&�v�^����mK�l[���R��������<E��ֽ1�i4=I���!��wf��Q�#T��%E�����4�U�CIDQ;�y��HBk��.%Ί� ���Fy����%��ufu��">��*pI:��\n`&�H�*�$j|��ߢ\?���䔩�ُ�c9�Z#�ſ]�d�h:7 ���&.y���� \}�7�����gj���e��̂CK0�)b:�j!3<b���;�}��N�����c�6��r�_�?'ciX�i�+OYW��Q�>jl(Uq���`җ��CH%�I�H)O7�Ǟ0������{��E�$��0���`��d�U��g�Gvi)���O�Ϗ�*aED�|�?����ñԈ�q:�*+ŸIZx�`'}/mY���[��V�9����-���9c:s���Y�&�=�	n.����r�Y����}}�(��r[s��AV9��*:#�UC�9��|��������1�H��j^(�0`���C�i��N��I�&���w�NΉ
!1�Q���J�κ*���V]����&�,R�����$�{X �wVS������w��s����N���G`^��[|I
�<�����򖤼��r>I���>ۯg�K��2�*]���p�Gȓ����vl�d�e��p14N�����������c����$�q=�
;�8d:NltD�dF�Tl���v;����ԇ�Y����q*Q����O=p��%�Ү���$w��u�~�_	��t�t+�����������kS������_���\��i>���B�m�°i������LU����5$
�l��3D1�IV��$��Ҿ�U"������F�C"�o?X' d���EO`��ƻ�]�*�b.�!&�-?���R�C#)Owr��P��KӤg?���Μ���Gn���H�~pV+>�)%Rk!1	�,�E���.�<�������h�����%�S�P�#\5��'�(a�;䒫X�j��D���j�yh85v�v���"S�Ko�og��&����QX�L8�O�w�r�å��A�@Z��<j/+G)�]��ngkv�{���{�3H����G���vW^Pɴ�d�m�W;���S��E%���^���:����c�d��h�Ƞ�Zw��Dhx߇���s�o���0+�7s�Vp���W������Y��r����̰�/Y���&�pp]�)PR�S�u�?k���.9��C�v�cdS�_z�+�H�rp�E����=�_���Ԃ��#N�m)b���%�g�`�Pv<åa-�e�M����`��'�!s�cJB���N��F��v<�=suC���\���Gw�L���q/�k�as��g͕�
�u���nw}P����� N's:�eۅ�}R/N�.�Dz�V#h�էܤB�d^˪�B��@��bK���]@�c��m���Q�
��Q{�k��(�A{!@o���E�K��cc����A��ϊ��CZƊi�#����)
x���x������-��\#F,���	��ǽ�3�48��9nrԸ]Q;K��Ħ"so��8�CT�嘸��_ d6 �x4���<Ɠ�gq�S�Z�B��\�뽠c�R���`����Q���-�n���o[$i�M�bF���>(%X ��0�v����rl}���m\=������i��:Hj&�f�/�T�v̺čo�a���h�����������m�u��>9ծ��#��~ˁE���S�V�!虶K����"�#��;�\۵���2��u��k���%˦R.Z��Sx<(�,������U�j�)��B���0I��HARb�V�ǫo����5b�l#�\�������7��DE���q�W)�ȆF9�lQ�z�O���O��T~�OV�����|�c�{QDE�jM��@N���M���� ͆/i����$sN��.l@��UӨXo1��k;R�;u��M3Ұ@�\��,}x��}p��+Y˹�y
��t���̊�A�(��(���Tϔ�Z�̒BB�6��A�'����������}�38̢�e��TU�ՂA(�=�@����@���u=
�aA�-X��+C���zeI�0(�	�K,Á�eq�0�a�7dlA^쏆r�,��C�-Lee��4��/��OJ��T	�`t�e|(+��o��[0g\�F�Z���^M�^����G
!9"2��[t?���n2����-�{:��e3���eL@�M\|��8茒D�`��U��;4�Y��Q.%}=T�>��r�HҦ�lkQ�g��o��C]�Kf�2H�q�)`�Ӄ�յ����	Aӥ��'��#�����>��E`e��Ev���%j����\m0D��T���	<O�p�����QaO[����LVB��KR�X�4rc���:T��i��x�=ٲΟ��cNf��L����`B{�xP�ts�q�x@�lH�_�1���u���z破�m�^B�����Kd�U��\���Gב�:Gd�ր�/�'��v�&#c���vF��YXB���+}��+�"�AoV�������&y�I�(�}&�YL���C#�xK▨ڔ:k�*!�b��X�V�x�Z��OP[Y�c���1"���ճ�)�P�Ԕ��&����ֽ���l�w�d���U:UFk�e�Hԡ�?��ԟ�#��o�*N���iq��hx�R���Q�I�:�JS{�m�/��5w�	�S�J�b���k#XaS��ʩ+BvӶs�c>�y�ɣm	��|��h���'�R��k�f���N��Ź�m�ٷv�[�H�ɞޱL�V"q6^׌�NT�:��ϣQy;����sq��]�p+u�2J��V��\x6p�PV��'	��a��ךp�گt���R*M]�B�%�O�{C!�^[�!H]{͈�����j��64�\�$�n=1_�����[PЦ�%ox>�]Ě%P;�7[K��Яf�0�4��eX�Ɏ2`l�"Ȕ"
�Y��J��	\=��.�f�\�qPϝ��~��n+^�B�X�f'��	�N�eB�ycXj~�GY�(�P z�W|f���$Ԗ^��*x4����2�W��@�f���S��M��q�2ލ�8��;d!�0yq%{�CYZ�W]ê"j�b�D�jyn��E�b�d�@���oZ�D��	�Rm��r���t}���Zw"s�p���s5��.,�J6��L���Vz�fE$4(�.8 ވ�7е�S���qi)_�����ߚ/.��M�/`5f_������޵0�S����@6P��a�P8�E@�	(�;���o+e*�خ�L-DXv���!Mi����׉��~ȗ0�B���=�( 8�S�0O�p���m���ֲ�u"rd�Q�Dq�h��� R�Ly�{m��y<�0j+����=�ui���S�+NCb���QL�t���QG���b%�!6-^�C4��t���ަ�tk���!�h�Rd�Z�lU��e�k"\��	��{��$_[5�v���K03Z�叓Ѳ���n:F �� �X�Oc~.^
{�k����-���
i����^9���l�����ϔc.q浕*񻷣��2�B�8�S����@~��Z�.0|�6�(>7e�?��<����˹���c���O��nܱ�̸��Nc� ߍ���j�/캖=�؋E���ܤ��q=fEŁ��_j{�7�8��c�q�bM��,�it�l�)QJt	%�1�{�k$��ğr�E#�1��3����7 ��E�X��
��� �6��J�x;ڀ�}�!��c���C����U�U�M�	�z�^Y�뤹7�+��_ F��pF�e�� V�G�`�5U"��:"�����d��]��C�Tl�93��۠��rc�����Qak�PQB�x����Nz�I�z��5��m�����u��S����[?����̖D�>F&%��Y�8�ra���+V�j(	�/,��mfL�"�ܰ�Gʤ��Pjs���!'����'�̨��x�r3�N�jB.��#��F�d�Q�b�ӣؘ�s3 G��Ǆ�U�Z=N3�̻�K.qmg��-��T+>�E��>^4IV��ԡ=+��P�S�z��aq��r���;O�@����D��z�bpx���#Lz��4{ao ���d�~�
 �:�e�C�gBq�l��ҋ��o���|M�8����c�t�L9Ǝ1T�Y1�5�W���䰚D�/"�-��eT��x������������(ϰ��>	�;��eZ��r����"B�ߥ�}�!��5|^T	�w�u��?�A���.�IMF|�i�2d��#�t0*?ٱ���XR"�`B"��/p��o�
V�n�A�j�1�hx�[����xaj�%)����7�z�#;��d�\����]l��ܢ;n�����1�=o��bz������b3�/�^Q�
� I����
I���^����$ҍ��A�tdV�5���S���(T΃�K�3P}e7�{3�h�z�6�䖜(�P{��B�7��3Np����\Y�Ś|}����~�p��~�D�����_�w":X��E��&P�k'��FLd��������Hd!\�_&i:{��<C�%�+������O��^������|��C�6Of�YK�:47.OA�?v� ���압z�E(��<�����ir(� �<%���Q[�4��O���N��{ҵ���ٍl(��i,y(����c�7�z���F��1o�s/#oP�����I)��^a���Xo3N���x�%�� ��Ü�����D�E�7D+�y� ����ҽ��~M�K]߭��^����L[A)�:`?�X���ͺ��e��D�m��!����6�NS��?��ȟȟ�ĴBn�ޱ�*Ć[	�]_X��6��oS��G�Qc��PiS_O��`�Q�>�<�{��""r��m���$_;�К����rm����r��G\o0.��߉~��0�d�c�;f�r{ڛqp��x8&I���!�і!��7	��f��38=��Ml�/ (=�~d6�:udP�T�vz�)����᪼�ʗ��b���JT�$rۓ�&�͏�qFz�r��dfRk$��̩�4�s��JN`&u���HP7���Ù��������~72�k��6K�4�ݩ��抴��RO�4=�SI�أ��F�y��Ag��M��K ���kɷo+tS���C�F|NT#v8B�+��!����	jMȉaZ9�����<�LK�#���a���� �П�_@���fkO���[��"����z���G�$��'������RY�G������z�|zȉZ�'��g��D˷�ZWԦ;��9"j�H����JH� �9�n7����jb���X,Q���NH��!bc*�-^嫍���4H��*��֨S/'B�j�i�@��E��*�^/_�'��_!-��|����^إ�H�J��y֫���m����;�8�H������o����wp�.h�P�y*g@$l��а]VD�LJv���3	X�Z�p��2���O�3s&h�����<>)yA1�ui�+]�zFw�@`�2]��g����2�/���6s���`^�ޘo�'NUN������sLQ;�\`��@��E?[����o�H� �}(�	�6�x\}p_?�Ԙj4qJcV��m-��Uo�fz{!��,*��o�'�>����s׺Da0�5	Q�B�NX�2E��%�L�(ƄK�%KdxׁX>�>'r1��/�"��ulzW9�M�-,�G��T?O^���,�n�(	w�
�����������Qy�^j�w(v�Xx$�dio�()M��5���D�9�8�����T�����m,ո�[��}�"���ީ��1� ց'��P��~yYt�C��ԟ[�no]��4�i;����;i���
/UJ�^H����aaPe/`U����G��I�h�R�ߟ��}g�1���	�A$v���v��&4SŢf�������"/�FO�<�ҹƆ�F���Z��t��$�Z�0ԠU�[��:h���%�P	����y=c}�m(�*��s*�n�5��=��H�ß�I��?�ݗ/�x���ݛw����E7qm~��Y��� (�Pi�~���ZM�[�_F'���$G0�xg�ZXັyWQ������GT�͚��Y"V_��^V,�Qm[��=���egF�h�L�2��zQ0�D�vx�Od+H��Ϥ0[��z�ba�u�����$N��RT^�qo���7���^�u�E�b�*/���Q��>��+�gF�L������n�V��-�D]i	��H_:���Ա�(��~�V�y����:i�l�$�wQB!�4k��`-��!	��>�0{5��Қm����俑��wϾ^���Y�D��{{d����҉�ҋ��p_q�����������>>��Lf��?y��4��轥�)�T|�g��	[��Y�1thr�,����o�l�C��7�)U��UP�,G�0ӉXG�ر<+��K��x�f�b�l�ϴ(�^*�2`-Ս�;Mw��&iF�T+��#GCpϼC�`��,�M,��y�Q�=�?a�w�A�o��>�:����AƏ�:Yt9����ߋ1ԁ${��B��{wG��]4)V;}���<?wQA�T3��ɡ)��~����َ�N��C��-�L��u^��e���T����v���@�C�x���[Խ�S�/�lG+ _�u	�>�]X{�ɷ�~���kY�ɀ��|:�2<̕*ZE�M(�\�*�-߭�[��	���sD�����%����`@q	M}ʤb *]J5+����R8�U�p{�i}�� 7��|�M'}`��yƾ���������s�^2kMgө��� 2]�h���6uk�<�_��BEq�l�[������s@XsЧ���{*͚(T�S�x=c@2�XKA,6�	-x$ô.@s1���T8�a1�8��?t`�Cլ�
<��������&#��b,^���t0zz*���q�<��Z�{x�����i̦�jb�Y�r4�m��a�<����H$ۉPǷ��6�ߍ�3�E���۩$��އrt������56*pD�xS����g�j�ؗ7����[�#Q���lW�Fy�%������Z6���Ġ3jW��	쿃S���/pwM��3-k������G"���L� e�P�!��:����3^�A�z;���������O�g�Ǟ��MlZ����b
�2�U}�`��:=,�*ąwQ����TY�*^�y{���?�*MMF��mL������#�*6r��54���7QkU4�)�6ׄ~9��$�5�&ʫ���~��+��}Eѻ�Ć�|��rO6��_��������d*n�b�v\P�m��}�P���MD���x����Vm���嶞��b���?����-cRA��+c+Ȓ�������1�̇iF�5$�����KR����5���&W�B�(EZ.Tu{hGeR\k���4��T ��O�k��`8x۳�*��e���V�p���HHu�
�F�eS�$y���(T��a(q�s)-F7������FD����&߶�D��T
GN޶)���:_`b��1���Zz:�l*o�G%"�[�'���Ou�Ns��\�I�M��[X���t�1�tv�u��ǵf��?�IJ툜7q�E<���ț�$JyQ���-��7O(�ʵu��|�6��d�%�6ją�*T���69فÐ�7�
0@�2a��%j������	%�+<��e%ĵ%g�<҆��x�-�Q�����s��.��o�d ���8Eh��&��~{�ג��D��E�����R��1�N�Y�ք�A���{�.�|SLbc�zEMI\v�1<��G/�� ��Ψ���al?u�|���d����H��?Tx���ۖ�tBC��8q ,��{��R��j�XtkC+�;��̩�r}hc9�_���Y� �0"_�i��3�LS���8����9O��RIMjI�ﲅ�Gc�0��r<H�w�]�&�X�h�$�ڌ�Z7܊�%����r���f�8�=���d�^���	t��qz~~LeĀݯ"
��\ F}a�n-�E~C1�mA��|�y����i�HQ�*`�K�+�H�=�r|�2���+��Z��31�>��T��DTY�4�E�Z �^�_�D�AL7���`��s:��k��a�PT��0��.����O-��ݔ�az)��u��?�×��{�;��u�9
q�)
6�ON���oWz[��aXM�(,hZ=�}uH�}`GizX���e7��\��æi�{?(HZ�ۆ�Q�?�Uf���{3�ը�[l3"Y*���'���D�H�)G��V�-`X �S���8�y�[cI�ol���Ib��o*
�'���{B��'N#dt2� ����!�?���A�LU�T͝ )�聗I�*�������($@�o:{OmK��!�L�\��I����_P5d��Ģ]��F���<k�f~`�;�L�=ѩ_"�������R_W\� ��t}�3���l Gw�ny@��:}�<��$��.)w�t��G��/wu*��LgBS�)���BH��2�(Xy�G�<ON���2-��A�?����σ������������05�����˒-ѿ5��DPR��oL8OQi�D0�n8��p�5f�j�E2�����>�+Ndr\o���������U��A7ݓi]��H��L?S��'�s���Cܵg��fLV���k�6�Vzb��AX�K*���-����7�,��+�v:�v���(.�|��Y�����m4k���Q��z�v�����}< �f�h!Y��%�C������na�y�ji��&l� �I!τ��3m5R���-�/:�
a�z��W��	�����ɛ����;��L�S"�a�wܳ��v����1�&vzޅ��JI�(�9|��1� ��D�FR����FC�������HE:��^�s_��]X��H��2�7Ľ��Ak�d����+i��C�>1�?�x�߿N9.�ֲ���l1�V,�p��M�z*E�Ȼc��K�cT��yG(���_Tbp�QK������f�+{5�J�7l�х�is-�c�+kl��F�ڜ�����u*@�5X� ����6�J~L� `-o�Ч����-d�-M����\��kӅ0��L��c��#�\M�=Gj��7����]�wp�F�����F �����@S�g~���P���Me"����e�C���)G�M�?���4�d�w��#�&	X�q8)T�|���p�`jBt�4��9���e�6~�S��e �;�>-V�[\j���c�,MM�� v�G��������4�;'�~�{���d���h_ �n�>���x{᳋ų�ofَ�?7��E/�
X-�Ԫ���a��H��fi�����M24�8��т�k�̈�Oq�:0��3%S��6Hޥ�o��&Е�8L���?�5�ܑ��ցP���s@U�{%�eM]f�4hoŗ�0�BأS�Wj����̌jd�]n!�V�V�@�d)�
��!~0K]g��P@�R�i�z ��<�t��pe���,:�E�'ͮ�W��0�tү�<��z�[��?}��H��m��[�#�X�'۾5�0m��of//����ʭtƽe}n���=1��<-���"wS�D p�]�\$|��$�b��;I(�����:=(k���8��4v^�z.�W%�Ǌ7�M�5��2�3�s�ޛ+]+�P�fM�Bug.*�2�̒��)Cc�|�!��?����I5`}CE~�K�w�
}s<��q��
�Z9䅜�aBux������&�b�&��mi:`fwΕe�G�d���C�+S~4���5���#y�)�Dz���]��H��xE���6#���e x����o�8��m0)
�)(�a�Ѹ���3���U;v
�i���!o��s�-���I>�_ r�L%�)ۓ�;p�^ZV����C�w�ol��e��<s R@ԮH(�ͱ�+� I�����!܏�����5;Z�l��/r��<iwz�qU�˼V���b]lv����~|��ɻɨڝ��P���ĥ�ғ�O��:6�Rh���˃��O(Z[z����L����^^&�XoO���y�aV��tN�msy���Fs�����_�h��7乁j��&�%�.�j��kIt�R�ˏ���@be~��[�+a�!����0��h��V���s6��` 0��sB�ΟQ�ZS^�	�М�������'�(2_���ϵ�~�{��OE]T*�aͫ�n��é�3D`��2%��V��6����"��Oqd����K�u�1lߘ�t�T턱=@I����֊�#��������n��C)�95�j6�աC!��dpoJ�$����䰟�(T�kv�]���"����4h�E?���[]�B�$�p	'��Ce����;���Z�2��G�	7(�������⽰D���R� �Ă*�75h ���'Dz!9"G�`%�Q��&��M"�P��=1�ĵZr���c����,A��Iޞ��	m:�D�%���he[ �]��K�_e`��.9�fǅ^��q�����1��(B'j�����P�I��)Ccg�@�	�6��$_K����'�X:�:��$Zƶ|����ƌ���e��:b��DBR;�@��X���F�����X��ڤ����]\ե4������1@�{�k���'�qG��zn��s����Gcr�OI��vP�����	��ʫ��&
'��$�� ��w��*b�߸�<� 9��Y��kS��t��Y]��|͎��+�`�OGV��gt����G~yy��q�T������#���,��F���-����mI%�NIr>�$��F� �﯄��J)M�b(*-Uuo�'-t�J-��G�UP�eRȖc��8 �U>���d-�OE����-���02�C�RYiv��Ж�V0`�Ƙ�0�wz9�6��PBJ�
V6�P�ե�Y�D�cWZ��C�Ʋ����`v��4��3z{���y��j���C�H�=vݰ]����dÖб�q(��Q�4����2T�	��Kv�t�f�̠6�b�;��7�ݘ$�7Ҋ'��]�W����:�Y�?��0r�z*��O��n;��&P���=p�	�*�kHUe�|����c��'K�fo��i6J���d/��E��4=q�iV���az�.��a։�1��y~��./�kL����h!�֒Z~p'R�3co�DeVl�M���,���YA;D������G���(���n��0��D��@rt��ք^�����`�Rʝ��=��&��a�^!�F�r>Æ��S�N;�KI���%�b��u`ˇ���!�_��N�U�#�ǌ.[�^i������'ۛ���hf�5��q����E�aF���!.�~c)9DgliEoIm�u�_i�@ȑTZ��H�6I�M"˟r���RiU9���Ka2�o;%7��ں~�6xӔ3zC
+�Hu
���{�z�_
�M;LEbd�Q�*�-������?���h_�`v�R�:c�S5�Ǹm���NTצ�q_bj5��8�==m�Rυ�4�~6G)�;|WR���Ml!^��?a���̗� ~T�0Ѧ�v1�Xڨ��o���ΎǇI	ߥBu�˩fA�$XB�)�bڳ=H:���TXB�<�M��;-u*�����f�!��D�2����)$��2\�����p҈>V�T_�����e�$k�č u�����˙ađ�:��A� ���r���s��U�5�8�\/}�0���������iW>���"q����1��O)�P���+!DLed�}�t�o�V���q���P�ˣ�StB������%��e��������'lo��ޤ�
J{'�`Y.F�[b�;��l��_���Gs�t;��8N��Bƀ�D���#�w�z��ϲ�_���9!�TOs�	��EB�CH��g� �w��\/R�)�| 7~l�t�h��`���ua��P��j�GV�����e��ihhl��{ZA-3n�B�cI����&�����#�Rn���c�V�$z�����[g��B[��,��\��~��Ĝ�\a��Y|�U�D0K�j������(B�lg�d�5�]����$��.ӣ�~=�������m��2�c�c�^��#�<���j6>T�)j!�18��ʩl]%��~��vO>�y:���~␺ˌ��o*~��^=O�X�K���$y7!f��=P����R�B�χ��mjfJ�Y�ej�b�O��U�M��a,t�����q��gO�˘3�: q'�؇$ѝ_�0Mጙ���QE��!fr�ꑡگ��m��;,p�5��c��&���P�1�'��y;Q:Q��b�(�������� >��b�����pA����
���I�Q
��-�1�L?�����u���oR�ck�2��2PY{�5�����o�9�rz��p^��
�|��)9��i�0�M[�};�?��cegPU����|���[�%��j�b�����v��:����1y?���୊��+�1������'�t�쯱~�0�C6�����g'�Ty.�8^�f�ŗ���q)-�0XLU\��l�t
���v��%t&zߏ�@Ĺu������ ��&IW�!���4L�S� a�7 Q���*��i����T�-��Q?����@�k��{00��&�p!��תּ���˃@��k��&q��?XM?�IQ��Ѱ��״2 �cY�ϧ(<:KΎ��-��#�wB�� �0> 
�[�,����'^"�������tm\>��9�dj�e�,�]��OP�Z3˽�,N���]uȏ�/ Ke�4¥�z#�S��F_|��mV�el��|ёIx�?e����~���31r�//��B&�Õ"����_����`�y�~�~9�a����`y���}�'��3 ��>H9�GR�oЉSwY�rj�@�����;P�g����,��T��֦��V�MK��rDګ��^�+��7��+�VE������'4JUQ�g�w�,�2�P���J��%� �y���FŎM���Zy�I����:�?M/ı�(�"ulOD��P,�=�St\���Q6R�/mP�l�Rں�5<�o\��|�x�4ktA�9�Jd&!Vɏ�bY/A@)_���﹩���;����2YɭK�/��Aض��@��K&��9Ar�bu���U�O4Z�\��汎C��<|Ju��ԗ���|�����*ԦR
�s��᭶^5h�����<_���q��E'ι0ىq���#f:����$~���i�>ϭ [hP�M�I�-A���>\��Z(��M��X��ی�}$�˿+dҪ��"i�Pe��9�^3-c��f� ��U�Y���5�����/�:Z��'x��\�ҭh�Y0t��[X�Q�\�����?6��x���	t$�螭�(�@'yTP�q�~J�U[���S�v~CĶ̆������ڰ� XEw�z�fde��Խ�)�����{�9�h��ň	
�F��������c $��?\����{����Dz��ɛ�h6g�<�)���*��R�&MPbh�J��������-�=�n����rr�G���KIx�8<��)���$��-�yM���a�d�����MH�mr�}���	��Ȓl֟Tk;h0���t�}�iP[�/c�4��B��(8���G媈��E��s�to�y��L���h�L�MXXG�59�iz�X� <Ý����i����^�=Q�պ��Y(����Dk�6l?���ީE#|t�|�<�n%�l�1��0#l���c��k���؈�m��Cq����1��1�|���hS!��%*�4�j�E
qy i��-9IY$��~�����=��XB��a�W��B:9�Ԕ&�2$e�(`���A��*a���7GU�g[��q<��@	�����e�����Ħ�,+�޵����1��佖� �"$�X8�Z8]������F��m&�e�]��]ɮ��W1��<��*�C_s^��ؠ[��������~[�g�uha�ѫ����3ܥ{'����w��uN���N�-;�>+'7Ỉ
��"ze� !��l2;o%�M�I����G8G�B��N��̢7y ?a���P�0�n��x�|+�Z�"�A����5܊zi���3@�����k����j�=P�+5Ш������f0����B��,�䂃~�N�u�F��G�����H�x�l�,������� ��?k�
�2)��0nS���;9y�������@�M�T���$Х]�[1^uZ�tză%Z/~�����\e����WJa�(~%�!FV�v����3�}��m�x�V���e��)ߏ�_�F�K�X��ז��	S4� }G2�o�L�:�r[��Xb�EA�Zp0�{��k�b˭k���6�E-C����p�,A;�-HsMr�)۳�H�z��g��_���BSb�k9�Vش�������By���W�C��%���q������m���ҟw��۶�R�UL' (��gp��]��c�S���fp�H`���n�K�����]M���[�5%��_�ԟ���Ϻ���wϊ��2v�P1݋lG�8<M�W��(��Z�EFb�����u �"��&�R��k���f�M$8�/���؂��z��HmSw�"�_ކ� � (��#n��geUO��7�Agu���	 ��~�����[
�<�SϸpĄ��ߥ�����ƃ������Σsr�_���CB�f="V?����C��$�!|��m� P����2�i{�R
�E�W�(_1�g�i�	 ��J~��@2�]�������-u �sdמ��BGV�gLҨ�R���jKZ�6�����I����HR�D�I.)P�5�Ջ��f�Qh̞gW
S��L���Si6�U�ԯ��]v��+�Qɘ���0�!���g)�ӯ��7���J�*D��-qcKʿ)�|w��{˼��=S�U�KA�E�i�k6Rtsrḫ�P�-���>�R�v����p ����]1(�!Ufn��e@k�dX�ex�(z���J��"~i�
������a������=h|�+�l���Ky�.�c�ݙ���A�~�l+ٷJ�Gc�%���w}ז%�C,��4Z�2ހ1�HR6:i��33�1JG�Y�=��N���1�R�٤�?;v����V�v�mL�YV�����ʐ��<@�6I>�1�L�E���b��P�?����uxna:�;�����٫�L�e�;�ylqwY�X
������\}g���L	Z��C�"We;1Tfĩ
����<|�Ư'�� ���� ϧ��g��Q�r�4����|�~��ϋ+3(���m��v�s������|�����S�R���������B�R_?Y>ׇ[�}"Xo���6�v�lqO(�P�g�� ?ezf�-D8��/�1]��~��ڿ(���֌�p%���E����+�I4�U(�m�����Є���:�e}�˹�z��5���[��P�r��<����^�l����1F��7.�h��#�0 2<N��X�\U����kV?�I~/�xðɓ�(F�*��an�t��P���aͽ��� �]x9�����	�4����E�/�p���b���Np�n]�P	c���$4R�Ԋ�K���c�����S��I1��thQ�3��LEj��@����	��I�0���iy,�WnL�݌2t�H���Cq+Ƣ��;����?�v�V���ޖDk��n頛��һH~���;�7�gZ�WO�c�S� [�1<��}s��z�qIg�z0C��A����h�r�%\��$@�8�F9̴�o>���@���,Si3��Ev{*����`j��8&�*t��E-T�T4s~�J�hEK 
��ssQZxL�W���"%�_��SQsT�y�enf���g�Ca�QJ[c'��D=PS�_�"������ko���|Zh�[�[jG��g4�O���rK;�
��D,�4����<=ѡ�0/*�t��)j�e�_�gΜ�H͏�MVxf�R���E�lH����eQF�� ��EaA3����}濼'n%'���\�*������!�!�	"nC��~^�L/�p�fU[���� 
z���dwbi��$z���o��u�������t|��5��ڡ�/w|�pw���h���{�0��ڗO+�5��\�'���SY7�^���-Yo�x�E�Pvr~.%���0��������������ϥj��l�\$a��Bf���GM�%/�;ڑ�Zc����ND�O�;��?�$�v.ݏc>f�݁၀��xK��e5*u���p�(e�0Z��,�aۍ�TV�BZ���L�@"F�<o��2�Of�(�bSi�^"S�Q�߆YM�V��!ѓ#*jIR���F	܃*�� ���g���<��t�zSl�_�@H�n�Z ���g}E<&�ۏ�����K�7�e�K쾔Q:҆R���tX&����yN�Id�S�ak/���?���C~C�='��b�}=��fxv\���<r�i�{o&�iuG�*�84mF��t�N���8Տ�Q2 *�d�)`���{���a�|V"6і� !�q��X,zC�!fk��C��wz��Ӻs��Ձu�Ջ��1b�W��M�a+�?,;)����<��V��㳡�-�:�1���Z����s*y���Ғa�� ��ر)}�8�N����f�Xʽ�xy�в�=6K����Ws�
dN��*>^qwxq� �F�C��Z�$��c��#��: o?-��{E�|X��\�2��}�ƥڨ�74�������&�p����7=��l�1��6<����o���`7��݌=4-FD''t�ng^��?���p���l &�����F�P�\_�:�.�����P�s��q����<*�S�3ib2��~�P�����{Vb±�/����A��S�	����a�Vp��|Y�J��|���y3���k��Z�Fq��k��C��T�Ф��|I��Y�+�a������Ϋ��N�|�z2�O�~b��N��|�Q��,Of��ɐ�°&G�x�5L鲄J)�w��TO�_�dqx��i�YWN0=���ve�#��#��GE򺐃BXŌ���T�\Vbz��!j��MJ5���IQ��4�rș�K
Z���a��ߢ_?�	�(�+X�
��Q���Y�p٪�إ�)�̝����[���QU��Rܛ^�v,L�0�j���'�D���2j����_�/�R�޷�Jn�ʿz��
��	�����"�p!�}$sΔG{[+�&�����S.S5j�EU��Ux�J�tr�F�7h�^_���HY$��n���yOJ���^�`+��3h�3%>���Z㞣Ãζ� ��@�.y0�.�W�|��.vֆѵ�t0�N���w9��b*����Sp� �g)I��i-��[�-R��G$���D<�E�؂�K5�Υ#֤M婆�-�Ek����������2#�����q.3veГ���(*�N��N=	��J'*�a�������i��L�r̿��hCu߄��[@���y?���$�]?+1��u55�bJ��?6v��6;�6[��m]i&��������~�U;bK�F��/+��,�J({�"��j�^n��H/L�X�
�_���/Nv�,���;��ρD���]뽐�)�h+ɢy�[�T�	޻�������w��q1��L��g)e(�Tc���؂f`�>,�#<ؿ�̾�y�ݢ0e5g��%�H8�JT����NV���[	DqΑ*�h>Y��=��ӇX���G�+��Uf�2�����0�3U2��ߠ�:�5��m#��J9��!k������x��^v���G0����zU���7σ�%>����@:]=��8�0-���.љ�\����"�*h���Ь,yغ��2��u$���w����S�B�m�$~�^K����>I�"��Z6钹�&@#G�6�:�y�1���MA��qQ�R���G�Z�'"3Bn~\�r�ݎ8~f���̕���a^�q�ﳷcjc�.p�
�SHVW��n��a��sՂ���qym�	��M�Y�2��
9Ƃ�q|����'�B	�yŨf�$L:L�:�L_+
�+�Mq���3Z����[	P�ѽZv@M����~���||���OYT]+D}*��$��kRl]���f�m��w%�����g��fJ���fR1?QK��M��I����w�\{܈�܋߃���˻ͦ`67�jz�+zA-���>����O\,zY�]x��!\�����]�F�#y���#.b�!J4C�~�R9P��n�*֣��_H�%�M80�N�`��e�%'Q���ل�3U��o��5*�ˋ	���3%m�K3/)�k���P��b���+�*��\�Q&*Z�3ʇ4�����kE~a��>��ʧy��s!�D��K���� �����H'�ڀ�֢8n�N������:��|޲�	k����b��O��F�W����4�sVw-<�­Og�|ZD����5�:�>
��58�)����jچ-��H\�?}�]X��*��\�K�ݽ��E'J��?���'�	3�!޳,�B�h�4ɼ�-�V��A�����7<��d��j��O7�@5:ڂ�>�nd��䵢���ϔ��>� ���k����yck��M�����r������ȥ�=T���C$^���'�]���� ��ݳ,"u?��XA�Ӧw�n��R��5��صWH��v�����Npc��0<���`�Y#��R	���x�liA3>�N��5CR��D��80r�to��z<��DU���c%-�=�2�qZ�J���	���u�v%�� � ?�\԰wPA9���Gd�.H�����!����`�}�0F��˿���;�5��^Ϩuв��z���H\�l���J�#^E���mQU���i.�!B���wAv�fL�4��Tτ��Cf��ސ)8�m#��ncu��w.nE��6 {��3����m��C��Ke�y�\Q�͉q��W�r+��9=�,�k�Ū�C���k/2� q�@��o��=�?���~.�GOC� 0��ev9������j���X�O��&W���[-wy��3zK���v������S�������%R��Л����PZ�3��=��2_��IX�\ٛ�XL����m\1�V������C&smi�Þ�o�5�w��R�4�ه����'�|\�Iiyb$��b��gȧ�`�c)�t�O�G��~�e�!� h!���Xhs�V���鷫/��.���nE����v��=���n� ���^�+YG�Uq{�Q�V��8��.�`l>a�h�L?e:jhQ���[d$�R�+�������#J�t��ո4)sbM0�.�۟�U� �?��D�AF��ȃl5�UR�OȾ�^���1hWi��X_k��5�_��;"�����`���� �o���~@���a��h��yS�<����g0���G�X��Q����~�`��� �s���z}}-r�NW�dF@��q�e�*_����\���P�E��,cʒs��'���uפ�t������{נ�oR�[p�|�3Ak�᷃��J:�ᾷ�vR�C{Q�Xd�`ٰw��'h6,�c�0���K땧�w3�>���H�+Q&�۝��z�ħ)��1=z���~��I��灊�2 Ir�5�)E&l'�O�=E�V���/UblԖe�8'�Z	�I�
]%Y G>�V<`/�?�~�V�e�����%�J�}������+���R0�:�3����x�_�X�A��@�+���)qs�tիK�#�(�M��0ʀ�O`�A���Wc��=�V��_^f�,+UW�t���O���`��죙�2��s	e�f��b�Y*S;<���u ���8��ݥI��O���~;v�y���C��
�*�L<2 ��{ٚȁ��/$�-� ��t���r\�>U>D�?�]��i��p����~P�8!��[�y�g'��iWj���P,vc����M�b@�#���ݠx���o;�ذP�C3�➘�9�'�p�$
�9�ǃE�����%O�/[�F��œ}�,���>��90{�d!/Q��f�%�d��.L)r,��B�D���r=���`���Q��u����� �5�5�b*z	3����|��|'�q���+|�\���͒�<�J�Y�z-}�Y�J$'�O"AGtt�B�R:������B
TH���}��0��o y���"0��`��m��~�q��`�E�/v�%�����]����ҹ�:�� ��j_�Q$i�F6�_J�mϩu|�|��m�ؚ�tZ��e+A	��VAN�'
x�o�'�R3��/��@�z֫�ٛ/�D�y̳�~�R<��
��0ʪ-��;�`�8�tq�;6ɥ��=~ҳ��u���/�f`"�1M���/�8惊�	��M>�YZ��X:���]*M�{��H�ʴ�^?�%�.iթ;P�im�����F�[����\�!J��܈��3L�*�,��-�QL�{RsϨ�!��2�7e�@�I��C��,Ђ0�B�o#�4��\�L%���оiYt��%6����P�A��~K�ШfO=o����6���Ҁ߫���?o��Y��M����ۖ
Ɔ�6CR���}Y��K�
?j?x���h�)9.3Z��j��K �f�c4\�?M��`Va�)va�)�~�K5�/�Fa�-����k1��.O�Գk������wy�B�K����:<tV�|��C���"9t4];9	�?�(D'#��t���a5�|���yGm�<B>��74�"�ބ>m2/,���'Їt&0��E ���ڞ\j��5����p�2FT��p@9mIK^U�-�K��B�+�	5����M�![����3���>j+�t�jN;i�?ϐ�P� ̪�B6eʠ�8�,�+p%kp��X1GĀ܈�ٰ	�,V+�1G@暴��i%��FD�n�D���$v�5�
��,P���ϝ�=
���Cz�����YR{�I��0Z�"�0���F���/�T����X�DvS�j���ЮΗbP���sZ�:@���6����k�zxA_�!���h`~1xpk7��K2M�=&��*�-*䯬�u�+�̿����|��d%œ*�W�rH�ke�N�U��
f��-�+���nR�Ly�Fe�:�J//�]~��ZΡ�����VE���J}"�be�)���,}��q/�#NN��=*��$�=.�G���C7�V�L�'�;� aM�)1������v���tNR�(}y����%*�ANG0�#lt#j���!"�a��V�N�s�a�̃�}u�`&�҆�e�~J�d�]�̆�JYn�2z�{�B���8�,]x����R�@��00my�0KeKtad?+3��vc+�l�-��e���-�n�sjro����s@� ʓ�������B� �"�%I�2�-"3�~���H@��_{Vp;�:i�e��L|��(��x�����M�%j�?�`��
���ϣ�"�E)����@;?�j����k	�Y��P�Rud)���/gh߃��FR�8���5='xŻ��G�/��"@,թ����B�sV��!�ԯ̻��n��e�K&�\�����38C�PFGrd54�(����<�d���ȏOzu�c?�d/�]���T�!�����˦�_�0�����쥕��:�G`.��]�q\�V����!/��r+�]�V�q�		�v���k�ECwsv�������,k�Ğ�t�J3*d�a9��d	��ݜ9���&���YƝ>Ş�p�N`���!���4:�N��I� -��ᧅfB�"�8�[�~.�Z��ʂ�$���p�b����1qrh�L�ײM'�VU*�6�On?�jZ�}D���P[�<�5��I�gV0ϕ�C)����7��q����-��Bo���pa���YS�|��;bXuD~A�#�XM�	�n���A�Pen�gF�H�Vn�J)K����z�.��Eb{����B�K���`ˋm��"��(�nW@��J��T�
#}mwE��Җ��G���o�Fb�=DM�P���?�P�2K~�:�NA�-b`�;8{m�������m[���9m:7Ku��ef��B��m�$���l����4(4!�Y���ō�5����&��>8i}�㞔Ր9�DUN��K���騀�}����ٲ����iG���|)&��Ӷ`"�ϱC_D{���>���l�uB���"H���<ݵd���S�	����v<�,���3:���-4yS{�+�r�����Li)6,��
;V��$4�ţ��u�"K��j�������~�M�)�_�������3i���(�N����|�W��)ç�"8��;I��(�P��z3�T�2���xK��B@�#b���2��l�F������jyi"��|��*J"�3�����u3�f3x��5p������3��_s����g�}�Y��.�G���h:��A��KEJт|�ý�$V׌�?�]Qp��z� V�ncC'�q#5�Un��_y�\;�i ��V[ƴo�����5����(Y�.�r"P��ۗ�7j��:�rTw~�Z���2U �.��5��Q�&��=@�����4z#M��f6ȗV�3h�wn�k���`�,�q-���OP��.� ����ְ��M�BHx\��$T�%��u�o~xj6�gWb'2�l.��;=���;�SBjy&��?�S�!	]JݙH8����� ;|\��h�rԕ�C���Ր�>�/�aG9�`pe��.�x��j�h#K����C�A�?� �p(Ղ}�������V��4��A�ֺ�o�F�H�
�1����*�՛c�����@��^'1)v��0"]����:���C�x���u84ҪzR�%tJ�nlSs~k�f≛�$�V��<J�,�ۈ���.Dp��Uy"����<�µb�H�ȳu��T̢C�,�r]�x/:��(�^n��t)hڶ�~�%~6_�O �zh��|v OK�3���	k;�B%��YT���MB֡܀O,l�I�7=98��OŘ�G���4�<넮@T�^�M��W6�N��h`��K�L?8��1���Br�D��`�7�j;D����䬈��T���\S �}�(�ڶ�Ė����/�F<�*��vi��>�]d�h9o����&$G���C�e6��s�i:�p��G�y��tv�+ߛ���`T~:J4�d�l��
���zT5'[�0�q��;�@,���+OuW^Ê���lպ���FU��|��Z]E1��'],;é���p��q�l�-k��! �DX�Q���/��x�����ir@���}^�F��3Ⱦ�CJ��(���>�PT���rK}�~�XlU�{���<��u�;��l{� �Y���p��^a�W,�^�N��-�ΰfF7xn4cͯ���ʌ�8�eC8�K��zi�Ư�3l���?��n~�'���8�#k��7��W�Ds�0n�r��9,rJ�e��q�d���\�c?�}��R�$�;�Z�F��ؕ��&���}� gxMpd؄Q��c�Zz��8)G%K�2���� ��� �߀��k{����C�=��%H�����!��J: �_�Q�')�oV_jߞ� ���k;��s�"�����-A��?K�:�ƈ�*�DW��MN-��������c���K�p1!�U�t��x�n��+	v�7m�^�?�oR�Q�ذ�ʴ�<L#�@eD7�n��vBL����.�.)��ZF8t�t�+=���j��҅�q�ax%"�6Ӥ)2+��b��z�4JЕ��F�Hj�l";�W92���&�\�i)�U¥�8�� 8d5*��F����?GE�A?h�8�k��E�.�7j����bA�Zd��-�����LF`�]|6F�;���-/�$^��ik�h2m���(sG��++Y1�}��?fOw�Aܪ�'�@��a��1<���&�T�z�LT%��v�9%(�z�c�� �H����P>*<Q�]Q�d�Q� fe~�p�4��iu��%pg5���{��E��t��\;G:�;�P�$�2R�G�iY@��k�� nWN���ll�U��?��w�m(x���=~r�䫏8F� �[;c��e*ŗ�\~qg췯@��9��w%XXVZp�|��VM-\�C4z 7ɐ��?h5��ԙ�r nFl�jf5l�o�"n�X�����u��%�P�]"�J~�r�V �l�é��v|Zc�T�3�����OP�j��u`7���Q�K1`w�k�M �W�������0[Ѓ6�b2{MP�8��9lY�F^�C.a���b
��љ���B~�~����}��R�'lH�FXN0G������\(ƿof�N{  h�Z��u~���0��m�}/�*�Q�U���-�e��Y�+���Qx7��XB�xX��-8Z7jV8��fT�ت/xJ���%��i˻c�����2�8���,cJRg��$,+���Q�
��A���0rof��Hh��W�5t�3�C�J�L�G�U��Xf}�=�PFn�l���H$s,�JfIGAF��%���S���v_��J�/�ЭZ�8�`}��'�B}��8�f����g�w+<_[��O}m=yQl�Mxˢ2N 8��J���(�9�*�+/HK�,i!y6�uBI5�o��ll�(>�R2���YxR*��4��4�0��6������G3?���1o���E���׃�R�G������(� 1>�>wG"VR��b ���a(}�D�K!��6h�sz���:�S�k�y�� ϨF��ǌ�VP���9�6�J|]n�Ed~�� >LRfs�����p+u7�y�x['�2�����55���oXw-n�wH�<1���ʶ�14n��
�����\RT�M��.	S1�y�vb�3mٳR.H(뜁+'~�h��^a���RRN��V<@��:+H
�	��u�
>�8�آQ�����Q�>�c�i���7T�(�ک�`7�q��"]��c��JUa+�6*������p��Q��w~C����t=���	|R�CLJ������5� M֡#���H?��-*�~ߚ��2�+e�m)Z�~ [M]9A����.�;T ȝrScdO&ng���\�.�߲V
���/�+C=_�����߭ݵS.�F_�D/q���/�Ŷ�4���4�Q!S�.��0�^�Wt���d��꒪]����v�{Nh���]Rim�-��w�Qp���$VvĄ�X��%�ԑ#��Fi�z2�;\��e�J�ߴ�B�M�f[�j���XO�W��|�f3e���΂O�@��o��X��l" A����Yw��%�ɪX$Y�ɨʓ���a��ˆ��%��<�,f'�L�f�9A��d�ƭ+�*$�mg�� �!�j?������� t8Q�d��S�%�!uH�xa)��;��k?6_e;��}VX���^U��k��2���e#sz��_A���Ǒ
�ݫ��顽�z�N�\�&ҷ��_܁{r�r�v� �@��"������d�A�Ő6���<��Wu4����S)�|p�Tʊ�\���0���j|���X����PX,\��е� �nR��Np�I�9�"rCYY%@Z�.���U��qZ��EI���RYf����/@��L�6@\�0`_�%�fw�j��H���]#��1��_�e:�������_ϐ���/4xB2|�B��=#����� N�OQ]��b���%ٝS��![r(��:����H��~��ф�K�Ͻ䟡�������ɍ�fc�JX�i���4�̕� �x� Q�@a��iK�r&��դ��I3���w�<�q��w�hB�9&[��+�s�F!�?����r��b���a�AC����;��,t�U�B�t؜����� I���hW������I����������B���1%W$t^W!/�t�בPW��8OV� ��b1�]��Y�����_~���ؗ;�+��v��ţX��h/��;C�R�=M� ���_����zQ�6`K8��r�uR5�~��Jw������؂!<����)��b�_�t<3q��h��۱���P�-�c.B�X<����}p��hd��:����p��m�C��@R�������!��Re#0�a_$�_��Րw��nE*c���0�u>K��I���V�5#ˮ����X! :��cb����P�����@	��<p�N�.�a �ͺ�T�
��T��񗶈o�4�l	՘��5��'�����mT�q�K������z�R���7\3��F�������+�e�	A2�=�Z�a��*ӏ^=�´�g�3�yeZ�\F��=���[��7�$ �[]�v�d�0�(��T��)⼴eC�sz��\���CdF$���琝��^|���#OM}F�4���u[�/��!��xB�I�0ho5�����;�d�m�m�w��Ns���؁���y$���2�+��j�W�{�8.}o��R���*����*��V���"Ϛ}�*8�:o�L�e�GYzfM�d���W�_��
&r.�h�.x��4q7�@�H���JYm���[m�(�Cm6��*z��Č����j����$���1��v猟~�Q���J~�J�L'��,:�I��}+`b@��F32� �Xc�q��K~*3c��e!��/�6V�a��B�?a��hJ����Fq���k.�"/��/5o�w�J6�KR�����4�������|�A��%�����ߡL�M�Q)js;���N���>:�0W<�膿W˔��ew��Vm�8�����}9H��=�2�"`�87����ⷵ�b/'�
�4��X�A-wP�+Z�����F��B4��P)���;_��%;:-���������2�b�C=`�˕(���7�z�q����]fB�][]T��w
�x��;ޟMr7�<�(["�']7��،�hvIW$�����ʐ]b���$��ϳE�/c]�q4㐃1I�$�:�f���b�#-�{����K4��;Q�Y��6�2����O��I���&m�e<�K���T%"�� J����w���aR�;iƩ������"�����r�A�ed��P� 5�0մ<��� Xę>@4&U&�{�r��T���5���[F����{�.��|-��K�ǐw������jM���n�u����|��>h�����7a�gX��G�(?�}����!�xF�����1�P�O��0�Ș�H�M��+j���~�J�J��l�z��a�:�N�2C�D.���o;#��^�i�:Я{�Q��5���i��
��i�>9m�5$a����������n�ՠ!�&�z�7'c�)y�fN��v(z��_hZ\l��"���(� �� �|K�aX��)��R9��*!68q���#�v6����I�}��~��昁��c7�"����sU�-��e?��AՉv3<�Mh�[(����JCUX;8Ke�B�~¥�����fB��K�k��]��媭�y��58��c� 1����l;F�� ��;�L�Q<��qi����ȼGO���{�����G�D�*�@��\��_T��$S��`�0�w�"	����}�u���+���H[��d�����k���b�Ӧ	��6��7I^��p�m��?�Ԍx�$	J�-�5��z!��܌�]��-`�p�,Z���#m�>�=C��"+����"\w�Л>�<�ڎ\s�gd�*&C��DH���g��qxT`v|[��J�a�
�@&34�o���M���/�������JI�e |�px�ãH�G7>�M/hd:�kd�$K�Q�� ��a�y�d	���*�.�F�r�,ѧ�BQ���R���=
�V`B0�T�̿*Y��Yg�j���1* Du��I;M}���i���"��q_�ަ_MMR�g��Yq?�����-$�2�&�kS�|�|��Γy-���Rd��hz�]~z�{c���7�يi�[��8��h{�#�!��{��R���Z=:!�čw�P@�{bREܡ��<��q������!9�W��ԖR�P�\�+zO	P�Q��`^ l|9��[��]��XYc�̛�:Sr�w�xo�TNv�pz�eq��ɦ>_9M���k/W~1��|�؇1�)�SPi�s�蜅K�]�#�F��2��׿?-�E̵v=����6�jT	w3Q=���\�&y�oI�~�.Ast�U3	�-�)�W��'�A���̟���.OB�dr�M�M��ǯ�Ë�_S���g ��Qo�,@�	�: Ry�N��������(�@'�]�)���=+B�84��t������da�g�v/�^��ωط��|�������|�;4A/Q�|�$
��l�5�w4�	��oyW�:�(6ѥ���!��L>? �;�$��dt��]��ẻ3��;��|��^��\��-e~H��Z�wA��7l�a���|�z��q�l�����(Q!V:�U�4��o����	$0�Y(��_�7Y$��[�5K|0a\�/�L�Hϝht�	s����=[�L$��_�����h8�y�g�֓���*��x}��a@�#���Y�Wq��{\kFk��{O��cw��0�K]{7F�g�g~���-��W�=�ޜ+����'���~Pf�0�Qg��%�A�.�U�� ޫx}���w9������ƃ���<������pAg�=�6-��^���� �X�i�B-3\�3�����_��6?p�3_A��J+��s_�`T7+K]���׻���=��1��,X�J�h�ܒ\)�DP?�*?���3���N�OFFFRGƑڸ���̬]'����5�5��4�+��~*��	0U؛���!Zo��v񊖲�;Ʀ��&E�O�2�5Π
�c�8VcC���c#L#�N�Nx�����8���}�@��ltݬn��/J��()E��{9@�R���z9��e5)1���8��+���O���=e0���$�}#�v1��.��P� 9]7I���
ha5�j�J&�:-@o��7�rI�B�Մ�{p�@д�;��/��?�/%���~B]8+��tJ��.7��S��\��jnf��u�D��Xg􂯚�f߱`�9>2�(�S�s���׫PX5:���-#����Su~���?#p��
�	��G?���<i���0��&W�>a�P1��)n-����26�CI�����㟼k#/��'S���7�������U�D~!�����8Ù�$�mYF�mZ/�W�b6`��b1�4;=�֚+��?V_8<�y�>`B���S��P���F���Zj�&�HI0|J�2hj��o���5uPJN3SV�!X��"�v�W��Y�?,����:��ZԊ�5�e/J�O/��[�v���_A��+�#��ԴO@s\}��DR�-�.0$=�}��y���)�ҏ���-�3/�NE�1�x^5���/�	S�<��B��g�V=��.QWv"��ǵ�3��NN[�����ei,hqI.M.ж(do�c8�W�9 �0���QGԀz,��U� �+U���"|�Mս�Jf��&C���i�%Xx�m��"[��3 i$m̳iR1����b&k
"�����`�����X�k}�x�yR�3E��8N�� rV�i�o��l�zm	����0�k����?3t� �%?l��|x�E��A2��V���J1�;�<eh�9����^Y_������mj�Mj� �+؅�̦M�$������y�6�f7)[���cP�	.�C�6�g���J,�݅e�����NWug�?�^�;Y��7|���hs�]$䄝�ڧ��P��G1�b%�`kܹ��Z]5ݨ���s�&�z�Y�1!K4�K��9��v�܏f��uF+Q��6�T1�l-^��yD���'�a����?+�g�,ԩ÷��GO����r�$:^�I;v!S5ò��+�q�����\��~�	����,��IX}�����+��Bk����IaɰJk��t;�"V�S�@�8�@]�E15R�0��D�Fߠ����5���*��z���ͳ%�.1���?ԁ����%GS�����M�;9������_�t�*�X�v�iء橩{xlز�6��u���c��z?+DE휥�D�9��3��|�9��ŵyߟ"1�E�p(׾K>қ<�.�k�
��{�)�'�Q僫,y^4��.�D���㦭�h���C���K8ЗѲ�����4�x,�W�N2u��M�����?C�P�]�h
��|%fv��[�/��t��aD�q'b�ĤϢ���:�/W����HmB��|�=Ҕ���WH����Ǆ��$���q+��iላ3�&�4��C)�+¿/��rU��,�Ǘ�����$�����V,��ZF�+�e#t�ŲeX��)-���9M~�#�h�%�����v�?A��c�fEe3T�� /;yf�K����^/{���5���o|�F۸Z���K� p;>��U-�t:W�G(~�x��t�*�$]��ە���
���١đmre~�Xh�r�Ot�6�X�V���^R��A��ܐ���|O�W�-ܙE·��54p��R�A\�L��e{���Wx�"mW����5��k4%���Fls&�Mu �I�U�Ev�4�'�|�����S�[PUv��]�3ן�T�����NZ��� ݸ���"�h0�� ��
'L8&��X~���8�:�'�`L�ڢ��G`Lwv���d`,�kܐ��A�͑^f�N�;-T�\�H_	8jZD��7��]tcx���@�	��q��O*�*zZC<p�InB��9h"�����c������x"��7V���'H�H9�>�	���0����'��ά7�w\�ɴ�Sr.�D�kLyS9�Q�z��l���4'tDǀ���,pN�xT��\a����b�`�"�:5zAl�.�5>d_��x�ٍaNu�	,p�k�N���QjԄѴX6^#���(T�]7C@����c?���ő�̇e��T�m"��K26�}ش]���`����Yr�ߌ�k�@w��n[#�6��fjA��l�	N�"W����8̬�%�Hٟ�D�i�J�6��^�;U;q���5cY�;i�M���}�2��T0q�@D��]�8b�����!d�i�M*��Jn��w?`pZ̝e7gV�OU��QR����tV�ů;ރ�b��H:�4�H#���|0��8K��Qσ�S�3�ſպ�y8�pJ��>�d��bX�.D�Q��J�=֎=���
-Bd���Ax?�MD��r��i����
����V��KJ�Nٮ6�B �N���{�H��h4�27��'�9M>��ݷ�z��4�oWF_��`�xRG�8�o��Go�ٍv���`�x����I�x�Ns%3�@߼�l�x�����+mw|�a��jv��g6�1��ޣD:�M��8m�NO��؊}f�V>����d�н�^'�b���:�H�I��7Qbt����d����qX�-yU�Oo��ᤡ����<S�^#h��[�ٓbP��矆�re�U��oVX��qC��TK�̞HtjR�e��L1!�R!i�?X^���L���`D�)��M*�]`Mz�H�ia����,�_f�¸�(*�K��"�@���UƅO�D _¼ 狛�}D�o4H��ñqV!Q>l����_�s7p��:sv1A?�Z�@a�6_�9��%�1'mhv���\�k�����1�q��*6�Ӟ���k#�s�J ^P��ب<f��1�B��rV�I��m(��e϶N�-�ǳa�%�����-�dϒ"�
�i�f���vO����B��9���a^�
��!!a��׈�6���p��d��-�D����T����G�C�g���2��R�A&k5||
�B�%_����d��	.��5�k�5A���}s6��x�Jv�Zv�)�Y�-&Ě�5l]�.B�9��Oi��=+�w�SF�L��G�3�$�[��G�k��lf4)��l�;&����K~��Jw����^��ܞ���[xtx���f�6q6��(���^��Ŏ����P�sF��2�S�y	Z��J"^���2�D\.�&]��/�0�RS��ЙF��Z�Ⳃ��^��,�(��E�� FA����vA�	a\��TB!ﾋPS��E6Y}�5ˊl��W�:��>����ҷӎM�,r�����m����69;�Z		���ߎ�̶�F���~�U2��Xv�y��TT�� ���W��mcv��$r,
Efd♉�5�9�6�}&��'4]gɛ����/��B�e����c�5S������-�|���X�lgؔ��&tɃ&ly�M5�L��J]) ��]�:PMp�e!�&�*��K��Lo��h��zAn^��
���jl�i3.w����=�w��u� q���{�pVj�t����p#q��O�>"���!ʣa��ײsWt��Yv���6��f>��=q6>��./phj6 �Q�tǁd�?f�R��9��F0h��H�ɾ���(���#�Xa�$�H�é���&_������
�Մ�pb���z�����q���Zݦ	`�`Z���x�Ŧ���0L��eö���K��9�2��յ�慷I�W���Q��=�#Hf\��3~����/D�N�Ix���]�"�>��Ê��y^�"7@�C�Okّ�l��6�!��OR�qJ	�������.�6c{<j��c�C&�d8��MM�S�b.�,��%a�Q�B�H�_�k�O~u� 9n f��Zß�Ί�/�q0۽CF�;o�}�u�20�Ϛ��:k�o�]�=>	��B�è�s-35)�a-%=�>[s(�O$� ��gR�廒����:�m���[Y|7�����
���a��㠥Y�;$��ܔ�;X4B��ۣU��\��;-Cj`�s�HpiԴ��b�9���'�_%�g��A�CH�R�N��1�ފ,'ib��
P㖧��I􂯖�c1ʧ�Ջ���l	ME_j$���3I����W�_���`Hp$���Q2�P���G$(1*�@=�pN����K��[�i�X��+�ޑ@�����3�B�<����W7�N�d�n�I��ހ��*9�;k&�Ժ�0ڇ2�1x�>};����;v�Tg�f�(�J��e��3US�M!Ml�J|1��	8�&��r�&��tp*/C�d.G��s� MG�ٻZ�B@�>r���w�h/�����ɒ_p�J�Rf�&r�\p;Z���&���鑱��;6�x`��	�����/�@Y��)��	.�H�?��m<Cq�(�֔��ދcF^�iT��:N���Y�%�p~p��ѳ����5�w��;>���k�Z��ېy�H�[����`.V�������MRzE��%�Y"��mtD����>.�H��uLX�#�M��?ҵENx�i�K��e��%��ωu�s}^����(4� ��o
�se�=��ꙓ�h
�5GlW�8Q�ɌID�6�.�3�����=q����I׿W�|�M�)�$��p4�'�:�H�U��ޮ.�ϭ
�sM����k�ޘ�@s5�[t:��2x�k��pJU�z�	�!@U��[�V�"D�~�lX�kb�����cs�`��݊PHԄu,��\Z�,��,�h�=Z�+!�a��}+�C�tW8�0L���yHc.@����z��Gï^∔#�OQ�-�M������F�>���\Z�i|'IvNI:���z�n,uⱰ���O��ł5��o4��>.��z���n1���;���Д�\���ϟl��U���Bn����m?�������=�A7.خr�_\�.Y��w}���ҍ����%���$��~�<O��J[)�#���<�4��K9��z�	��:��t�_ƾ#V�Y�r�	$wQ�[f �FM�Y�yD�{K<i���Z���eG��l�Y3@3�
~~��~+�4]x�G#C�#{]��ũ��K!&}����>t�R8cIH������,��D��@�a�V�HhԗPe;�;�H��x?�<� Ȣ��قx-I>���z*혟�X(�P)�l7I$dM#|��%��՝n�iX+G f�F�<v�};�����0}�\x��>��J,�q�tz'�ۭ��? �_�n�	��ߝ�Ҍ�]�e�p�F�n��]���t/��ƋlILN`���v�*�o�G��T�QÊEAƊ��$�u��{���Q��P	Z��5��.2��%?�	E��d���C�v3��y�`�@1V��"�kf�$c����O*ŕ	S�[_�1
��k\x�u�û��m�)rL����v�:�}���=��#��GT�4���o7ˆ�~ wB���i1�x!]��<W)�?��w�X?;/��'�I��<��s�����j�rd��k=�,=2�܃�PZ#Sx�s��"���b�~�Cg +l���ѐ�R�4{|ͼp���ܯ5�>���������D����Ň���}������~��`�]��,�}�����HO������lr��/��hWHz�-���h���B=ڻYV�^�S;��ۊ���2�y$7��@��)���`�Y�d)�/4h����rԨ�^���,�L� ��.{x�؁���$+%������ ��=x�X'�o���G��h���R�#M;3��bf�b��.�O���b{l����~�I�)*ɫq�GEI6���e�(��x�J�>A���̄L��i��U	��܏g��s+��q	e�f��< ?V���T�͛˱_��3��<�2L,*F�#F\q��D���K�9��@cI��0��l%#Svnԝ�D��EGC��y� Y�\
���?�C�A�~IԲ�����J�� o��_��<N��S�õ��)%	����+B��6s���@hHWq@o���M�� Gt��6>JÕw��N 8x�ȥYmWY~�٤�i��ee�W�E�]IиE:/T��T��]R²%��I"ݺ���3�ܭ�%�L��|M	�M`M�G"W���s�{S����k��ߏ�;}�$7�8�~�+��wz]v�K8�(��MB�����`A�B�w$�vT�	6Hc�I�=t��A�'��Yb
���R]1�@��Bd��<�ȁf�sG(	���������K�2A���NZ�G>6]�:r��������%R5��v,��>������$�ێI��Ns(�O�@͈�u��8�
�h&,�ё�	$ 
�lW/�t̔*�]STr����yӪ�.KJzq��:�?�r���w��Y$���I� _,��k��})5)�1k+-f;�c��+�ɼ�0���`�B��+ܙ��
#I���t�G&���q�u��٧:]��l��1':�f5s��Qx1Q]���T�=��Q�,8:d�X7�%p-�E�^1	@�~��|O��L��iD22�z�� Y��eE6�b�W����1�ro�Ъ��z���S`}H!ӂ0�ow��2�xk,�޲�{+�����~�sL:lX��f�œF�],A3��X���m���t��.W�)0{��ʪo���G�����o�A��%�&9cZ�us��Jz8�5��(��Oj�2����w��]��[Jߏ�"�$y��+�ƹhͱ%t ��ZH?1p�54\�����ӒD76rv.u�/z1Q����x�v{���an�MP��L����1�1`d���#[D.�����:N�n�Y"�Qb���l���sz&JSIs��M���\B���5(�h?5%�:B4�v2�	��(=X�*�,���`,\�����\��G��b��nۏy�ӽ͢�ܬ/�\���E��SX�<6��i��}W�+�8����b��Sc�Y���}2�)�@��>AKH��)��˘�y%]������( �,�N��g���dt��ɰ����\Mג��2��]�~����X��S5�t��ӟ��~pױ�=���I��o��u�7����+'4�v���l(s��C���jC�5��6�XQ�"m��S|�ϥƚ܂�F�`�8��P�}��m�f��k9�A����\�s�@;��@V���^�t�F�5W��9�����g�$�T~)��\�h(�W��T����0k��'�u,���s@u�n�H�"��%<UQ8-�&��[����t%�7�%�cI�H#VF����&�q\���U,h[`��]i���+�Po~�����dhB֚*�i��/*�G`?m�Vk6Ζ�W~���팶�I�ͱ��
p��'/���B;���_��O��Vd����o��;Em���)φ�>`�����
�
li�55�K��b��.X��:sWdHg���r1��V���[��b�r�'lc�${.��f�|�K}��R<�+����.RX}j��jf�ua�|��X�(���p�m�p&~ۮ
�W2��yX3>f����mjG�w�|�`��K��x�%~��\&.��t�;>�.���W�W"s�_2����J��� �+PT3};����j���:��RG3 �˹�i7�A�{vw���-���U�����먠p�U��6��>�!�N��" �#���yoH}ˏ�P����>�߄ƶ=p�l3��ybS����nx;�0���e�W�F�d����k�27���di�F���5	�!�s����P�>f�73=����t�pa���R�R�٤�k�+�J��Jީ���I�gCe�_���}�},�Wa�ǌE���
��Oo��P�,��AKV�-xg�%����a_t0�F��{T�!��lC�,�����b�]��_��"k�ۘl��(�����ՙ=8k+O��v:�q����}\}�_��Ķ-K-�3��$�so�`��@E\ *s1�:@f������v��D�:z]�*xʶ���K��1�-�W�[Mi�V�߶8}�K�B�r���tl�4�h^��	�G̊��hi�������K�| 1��FS�jvi��e�\� XUm����*��d��\?�i�F8���3���]R����ꢗ��Bs�3c����@��!"�5�}O{�7.�+�H��
ˆ�b�	aA�w��o������|ǂ����\�e���v(v�t>�D,�j���(,�0�Uy�r��(�M��9� 
4��d�l�y��x#��3x�l�l.��D���ŷ^9��?�m��$�@�"�¯k�o�%!���g�G<ڟ��*=MQ|1�UŨ8 ^"L0��#�N�=O��o',k�̰���'G�.W���>�AjOUX"Svo����������C�����{g�"�ag'�y�H����zЉam������ڇ����fX2X�>B��k��_�K6�=����mÓ�	>!:�*n��:�Ֆ��<2�]�G�JJ�6���?�ߒ0�@)P�Y��������Vm�d�I���ov*���}Q6V���
J�))��|��߼��>?�n�M��ҷ�1kI�+����������-0Cz��|S-	��Cg��O��$�+�i��p4?�?�D��]�V�I^�Q���`vg�S6^��������#��/��?ݻ���D�%�`@�GEbf�o;�!�;�^V?��"Q��M?wB����vq�3���4A���Uԅ��y\���-�d��)ɟ\�R�[h�q s8;?l!aH-�cxhyam\G���|��'d\�Sh��E�8��d�ln��׫C6�B�y��;7^�r��a=�*��ꠏ�@9�~�4՞�.`���Up	.����d7���0�(JͻDf��X��t��,��ߠ��b�0�ܹT;@��ᝌ���Ci1\��� }Da���)�2� 1#2�+4�p�0�٬����\Ś��:Oo��0�a	�q�!>F��jnu!��]�E`'�"c�1_O�5<�w3�T �8M��z�l43Q�ӿL��t�\�7�C��V��	6%T��A5ʽ]��?k��L�k��G���L�1�A��A�����ѣ �_`\��㽈Sp���A��Zb���əy�k~i3���p�/�|�']�b	,,>���hu>+<sE �����M������=�E��Y�ĉ*j��9�&Df�`�%������Cί�Q�G�)USXm�4?oS�ɲ����ԍ��3��K����W��tW�ٴD�ҥ9�� k�w��F�B��b��q|�rѝ7��YU���D��Ϊ������+1@l_ ����6.]��hᇆ�0����u��6����d��Y�Cˇd�/����X������#{�w�Yl+��#���.���z3`w��O�����&���јu=u��`� �"����(d(�E� �θ�*��y�T;0�<�F�~��'U(Q��	A��Z��$n��J�\���IlJKΠ�ӵ��j��qp��u�s��$N�!��@�XY4j`A��2�<������k:ep����+~߯�H6zjw�(,'^��� �B�ի'������ z\B5l����~Ԧ}O³r�8t����)c
f�M��-�Ḷ��i~��q�l�9@6.�kiṬ���a�T�m�Apx`�4)M�۞����|���?�TʟυL�1?�K6Pa��MC�f������w6\̭D��M��]�w4������2�Dc ���E���aK�Uf[�|-/d^g%�&\O]H�8��O�ͨQ��d)�K�]�#�V4�Oa��^��{�fU�Tйx~U���4,:B���D�i9ӌJ��5M((Ç�D���R��c�!a�J��c�V��"���]x�U�|C5\MX,��RFi��c���أϙ]K��������1{�$5Yޝ�\�el�h��V7*�F�w�K��퐕�Qͤ�Y�q�U�M�^1������ax
�w��X �dh�N�Bd�~8�T��EUq�-_��Xi���\�#]�[D1��1U���W�\���a݇��%�n:Shc�Kl?t�ήp1+r�������~U�}�]2:z^H�T>h�c>^�;�Vn�md��hO��\������p�,�����P���-�4w�o��'�����_��@��l�/)�4s$uL��-�E�J�g4}@@W�z0�L�]~���LuS�:4,B��~.���2)�)B>�b�
/�D-gM��0sD�M��	����ݕbm�|��[�¯$x&�U��i� r����N#eP��4/�ϕ}������)|}�Q�a]DΤi;�N.v%�ݸv��=`�\����gӸN���Io��&�h��7�"O�y����io�������XXO����	���'&2��\"�<�5�P�kծR��Z��_�B�;s�Ć�2=�2#�ި�xu�@����/ү�������eVĹ�)=0��M��	NF��v}���_͍� �����.:H"<s����k#�0�;��h�� �.� hJvH87.w>�����4��0ܹ�D �2G�
r,?�7LM-h 0��Z����؁)3&�F���Z���f��G��Il
O����1���r���E-iZ�G�TG��@Ϫ�(w�+��:�k��XZ0�py��I�w�Q��,��p��O(5j-�g+��]_�{O��J���㦝5@+k�|���iv+���4_�ߦ�K�ew�h�3�V �����?��J7����-��Hd])P=��%��QFPD�%�_���Q*�X�L'i��i�&�v�1�11����N����	�� vXa����Vc��a���&L;��=V+mZ���?�&�΃��	�{��#�	V�H}�Z�S\\���.|�Οǹ'�t�hQzb�P��bn�"^X�}� �N��1� �+'f�U�eJ+�ұ������poho�&��r�h��v
�����r��n�a���"�{R�þ�Rq�B��'Ġ7��a)B��-�T�VO����u@�g�%���j�׌�y�����������'�����uj��T���+���������r���,�٘�����+�Tc=�d��w��O�؝?'�\]���������d����[(nkNÀ�s��~H�wl��N����-p��\@e:~M�k��d/p�ǭ8�ֽq�Y&�к�����U�u���2��z�x;��������P�T��HVm�HuAS�����
����E���Q[��9d�zoy���1�4'7ϖ_�K�Z���I��~D2a�h$v?�cw�;J�� ���|J��*܊�F$�����7�A����$e:+^������:+�s7>�	@�i%M��=lHӚz�-M�4�:�مy��X��Cϲ�BLHSMZ[��.=?����ЖK�l[G@��ƞ�e�Y��M��/:��Oʕ���}�Q(C�qou�c��{����i�.�I(Y:�r,ϒ�6M��-��I����2Z�� 4uڰ6L��\�\�z���(ۖT�m��{�̏.쵈ٗ�%.)V��Y�vżQ8*wʛ���Dq���ݽ������x���,Uu���s�a�n�쥰s>k���`(���ؖ�*/�3�Ҹ������,@�+\����tW�=�b��B«�V[꿹<�t�݅m���S��L����k��ȯ<`�o��3��b\�u$����Sd�$.W5��%N^%��b��	c���P��(p�
���|��X�"XN�ژ'5��.��E���r�V�K'��NP�G5��L��I@}ښ/:�$Ng"@z_>�a���gp#�E65�4dvr�=�8���0*�;���'h����|�P�4x�������N輫N���5����� �E�=A�V.���V��i�(~@�-F�O7�mT�ט�-�G�Ă�0��2PW`Fj-O͆���V�e��z�K""h$�
�7��װBG��Q��N�/n|����dZ/ �o��XE���fE˧�#;M/��9�i�0��^�1��n�R��̀�0!e8��u��\|�4+ÔC��k���h�V�yd[e*D'm�N2x��j�j�v�5_O�Q����� ʏ��e�)r�,�E��'�4�r"(wC.�*$��`�p�g���B`wA..(���"M^@�V-e7b�[��;J_u��x��u<�#SٞzE���`\�&k%�di̖�i�ϝ��}���W�ne=��
8�{6������͹�ʘ��H� #����qԲ-r;w�W�tU����I�6MNs��s���ߖ�����[�%!i3�¨1TAm����Z{Y����2	�7�Xq-5�A�� DB{�B������6 n�e�� �
�v ��ҷ��-:H*PDO�X��=(y�6=SX���w��s�#�\�_�R��b�ڇ�v*^��*f1�N���;α�K�Oa!q�:*�DS��M����ն����`䲖�f��X�k�,m��À��a:�kpY:kw*DePس��l����g�{cga�d��6��T�!�4����]��R�Ѱ�3K˘ЭK��9�GXj�XV<�W��$zLi��K"D���t#׾w(4��i�h.lC#���GLK���{��^c�����(
f�=[�秹b7�	EKO�sf�U�h(=~SВ,n6v�7��(<��L�` ۃ���pj���]�t��R.�Ct�@���p��~�c`~�]ͪ~+���(���K��V8�K?�C$�+}�(�/Yz'��V����v�a�8�1/�~q%�}E�^(�v�����F�&�lyrZ�X+|S��59U����Qh�^E���%Ы�I�IK�%�2;h��^6�B���)=�����O�r繗���o�� qvvV)|X�s���'�������-��[���d�Si�[O��;�mC��r����}l�'q�#F6��%��� ����t�,�@�ͦ<4w�/PG�������r�F���0Ɨ���F��L7N>�����P~B�wnؒ`:��x�mb��2���M�q�s�
H���T�� ��*�m̰��9rf�-)�J(`�o�'K��H�x�͌��t�-@���c�����[����1tpޫt8��%�mP(�D���%)�*O<�*뗚�+XaR\v^�xD�˲�d��	7����ٻ�˶���V����k��X��w
)����7�w�t&���&��3��%��һT�=E�-@t�!�.�rO�Tm�4�����6`\�1���Ԯ�V싖���̌zH
:�]�係xq���X H�J����r(�Bo�`�5�*�}���Z��"��|(0�R���Պ+Yk�O�ԧ����n
2I�U�aj����� G��I���ExJ���	T��ė�XLCD%@�m�l+ u�g^n��C��_fY�2�5^���T���[��#�ќ�H��x�e��&<b-����djfy߮���s�ް7�r��p�l�.L��l����7 ��(�*}i���AB�e��tB��t��54�@rK�S/��A�X;���0�l���)^�t��O�\���S,KKrҙmS��SN�1���3����v��8�J&�j?ꛯ���0�	)Z�꿌 Sȳ�[�
 ��J\e��f7�"�J���_a�&E	�,�U�b����#����H�'�:�:����8��憠5����0�8
Z���Pd�k�f���is�0ұ��<��T�*�.��<
��'����5�K5\��R4d�6��х,�ǝ���A�o�t��ɬ]>
$��7���|�J(c�i*��_��x����&��G�A�5w�r ^��#�+�¾�0{Z���|	���j���#ڠ'f!�]��t˜9��ln�Z
��0���9-����`�WQ�L�-_N�0!��u�	�3��]�X�a��6vMhڜ��C�eYv?5�}���ނ�y,�ѭޥ6�4����Oq0x]���Ԓ6%r�^�������_� ���-��6������
?z������C�,J�?V-z�u�AG�\Ԯ����:���KY�������U��c
x��/�T����+	ڥ�Y���)�ը�烒�X��Ws�����2O�����X��B�ϟ���ZOFs���.�dL�u)�TJ��h�g�� J;yV��S���Hr�E,�kg>�|��OƂ�eo�v�EuA��Qx���R�N_��C�5�S%���/~=��=`�D��f���ux�Ψ`��NM����X�u�í5(�.,� j�Cj�(YՋL"��k�w_ jV莮���pF��i-�X7�[sC�>B]��-�ۧ��� F��,�>ׄ^=
�T=[C=1�@�h̸��0�gރ�΁���$�c�FXp�����2-��6f�;t�����[�4g�y'6��z-7������)���!����҄lA���e_0��hQ�bq��D>[�S���7?��<5���DkQ�]}U����ւ-�i,���f"��Dޔ	(Xf����+,{�W����+ V%Y��Jg��u�*��O�([����&��� ��ѫ�E۹�u�,:�vǾd�kUI�~�Fł�}y1x�^5,NX�V��b�Q+�l[Ra�Z^�V3�y̱�Ps)�Q��g��E��]���U�Rz�+0���Ò�\T��H^��n|�ƕ���W�%����]������Ϣu�"��L�}%�S0jW��R��ps����q����G��"t�����a����d��]������Ds?o6�G����1F��F�u�nkJ�EQ���5�C�h-�o������9�Oc��?�ֽM��'�4�O��,־P~�3��x���J����� f䟋qZN�`Y-�6��v�b�IW�O'*]��c�8���W��'4
�e���ʛ����I�&�VA�P�ƿc���_�B�b�у�&Z|	��ސ����h��֒�A��*K���f�-�a�Ό��B�ᴰ0�M��>4��(&�����"zGt�f�⑻��"�mL��e8�NwPA_n)Miq�Rb���Yo;a�f8>�>�btq���ճ�o�{��y:�`L���IW�:�I�wφl����D�p�H?�Y6��I��4k�L7��w�3eNc�f.ౘET}�Q.`��d~�88��o���)4""�s]����{��@��נ����v_�m���#����������:��:府�G���'�n�Jh@ro��1���jJ8RA
(L�[�Kg��l1�����,��wb�p��ɯk�uiӻKp����X��@|� 3 ��]Qܑ!�Д���7�A�����A�bfR�n*��<���i��8������^j=�p@�^ ֕Q����@�1*b��g�x�ۖ/��L���Ls��T�˷cʝ.вCvi�]� P �l��_�E���h.�^�[>M��[Ѿ��.�7 �B��t-c�m��3���z7sd�5s���"%�A���_����e���ɥ����-_���$�n�,�.]V�z�ҟ���<�E��I�B�+R��B�u�on q��̿�-X'�>#�����ʉry"�n�����,l�*0>�w*�� ݋e��{���4�<%�uR�ہ�͌�cD�!��|���'eitU@��fmF�`��#��d�|E(T5�.�����
akP�x�53s@��p�q^X�t�p?��@,������Q�"����݊��ؐ���q�~�Ј����W�X�{Y+��K�j��T��6��� ��8���a���K_ȟM��^k���T��"�x8��j���`��P	2��e�	g��6��%��`)J��s���c�b��&�R ��I4�`�I�i�vo�T�Y��%����]���!B`��r~9�^m����g�
�j p���1��uX�o-���V��Ka9W�׹&�qD�$w�_Eg���-o��ײ��@�k��*@�~�w����
>�Q�?����^ukfxĦK�M�nX���qJn�����`"+�Cвv_'�C����a�_ZBZV��C���fe�,��W�Y�4���@iR:�{BG엶Y���ɾCn�Y�i,s��z+ A��?��x���(��鿚����L�;�CB���w�;}���c>���8�c�+.���������R�m5�� 5Iw�@ܒkB�q��e`N�5y�{By���+����"�e��B���̿�f�WG��붇��#	�?�h�K-NQZ��3�^�Sх�߮T:5��P=
���l����~��{��{x)̈́υ��/�'��ϠqE�c�ڶ�r�T}��4:k���Ђ�e]E�NM;A�F�zZ��&2:^d}��Sѹ8hpȃ�Q%���:�M��C�p�~ԏ�N�o}rF�(Ô�L[?��2W�d�u|;������{��ek���n@㗆��_�&�ρ�Y��o�[;��^gD�����{�I�c���������2-���`��E�+_3����t�1&&A<i�uP��L^�o$��i-����ڡ���ǘX5�8�?Z��X�"���$įڪ��9�`��-��7����{y��.O�:YvX�R�jЃn���5��=��\	�Y8I�rQ�Ũ@;�-�w��?���,��S��	zp7tQ@�`e��~OjBO�z"%���ǳ��_i��������p�Ƥ��X^��;���>��'BJ��o�~��\�9�~��+֋�)�&!{��8P����M�;���}g\)����Ө2��9�:ai���uK��O4�PZ�^��i����߼R�,y�����zD�0h���~�ZB��� �_X9k�}�k.��+n��e(�̓������8\���V �bv��&��S��$|r��v��=��)�����l��8A|�t&�Mߍ-1����0C��_�t��o����	l-�̏�44�X�B�)�������Ym�
���M�{�v9��`{EߨD����4�sp�{�:x��O^Q��-M
��j�t��*|�F��f�OF�]�i��xr��uI2�pT�,CG���L\�-�V�P��
	SE[�T�H �ALV"�4댳Ȏ���LrN6�q�\< q�7�KbE�ީ�I�y쉞������'~�����v�畏�	�׈Wq0����*SițOĞ*���5;���W�fL�[iLX-�����ّ/�Q ��g0-��`o�l�g�;J�� �޿Evx��U�_�g#2�xs��gu��֠���R��E�:�*�zyv8�nP�Se���=�<�*7�^�6���#�js�@��1+J1#��_��J���]��9
��� ��J=-9��p�����T����|�JH��A~� ��������Ё4�"��p��!C��m'����%L�x0)H�K-i>�fc�3tC ��t�7+ˈ4��U���ҍkOCw��-(5��I<�����Rd��q=��]���~�#o7��i|��_滸��6��D��ڍ��V/��<Di�=?^�t����0�d�¨�WuGG=:�a��i�xĝבs�8,f[�;�h�u$��%`[���k�r��z�B�c�5hX��C��I�aρ=�\��t�=x`�9�������6��<mR�c�_8`l�s3��^G�@LIE�T��r+Xy���T=O���4@����nsi���1=���pc�69�e��Z��e����0�s��6���7��̫Jט���w�U��Y���_U�`,�<�w]�_�:Z����Cu¼� �e�S�;�d�˧�3`\���
i�%I}�Y����P�
�t�x�D�^���2%���b,��ňF�KF�I�E\��'�6@�M~}Jv���[�]�z��v��A�JQ�KeC߸I�3�5����e<`�t9�b��n<�����T�loC�5!�eګ�@��f���N6�=˄ Xx�߈3)�%2$"c�c_Ћ���/���RU
6�f,��z�Ȭ.���0�3O/�B�_r�`L8nH�{&�A���(�M!�f�fo�H�F�&s�X�2��9^�S�*�t1�_�u�7������[��7��Oa��
����<�Mm*���-�Q�P�� <�2f���gͱa�#D �14$���Of�
Y��H�`��i�;���ҎfY՝�1$N'|Ma�'#���=��׷���uXi�M�Cu�`8>�J�N-��֫����m�7�e�'��lu�֛�]Ǻ�����,XXe�B�S�~��)"�Av��b7�J��=�,�	�̱����N��M�'��m>������m�!���9�w�{�#G��p�{��zY� E��8{�Υ��Y	]{[�G���g������a�-"B����֧V��/� �����4���
}�I
�>�S�,���k����{a������X��w����J�@f)"�l��&w/�~f��x��/�NS27�`� ����I�6{� E�?y�D��B�S�+R��6��L�-�Wf�A$[n0,��]�]�#���=Ͳz�M���@8y�ը������*be�<]�ś���Z��k��oz��ޜ<����7�U��K9���i����_Y4�@�~�g�z�=F�)���i�C׳����1e�}�ƍ­R�}�D�E=	� �b�����/ӏC5��tCh�ж4�(���;�Ih�6ï�:���V��pQ��c�X3N�,��i�:8Ŕ�E��zڤ
	�(�x�s��՟��'Z���]T�o�a9��W2rNܙn y:��1�a�[o�l���<�w'�_�.+;�����w��{�ك��m���o:�>�3t=�
j�%�����,]�B)�rQ�6xd��!}։!>t�/�+?>,hڙ���r�\E���O�?�jEs?M��5N�z�ƫ���?��r�-���fz�;s@7&;�](A�0�8�t-�|r��x*0,��m���܊��"[���B�:�Dq��/~-��>U�h�TO��D���]g����.(6�{O[��,�b5M /� �� A�8�"H���aB�Y�i��5)�?����ؖCc�`�x.����s�)i{��P�������5BB7g�\A�b�Li5�'$� �9J]1���T�~ � ��GJ��ڟ�h2Q\���F {�_F��$��f����Y���[���ٌw�եt�����0�����z@�Mz�"�ԩ�M���gq����XX�<3ձ�B	����i_FQL|�bz�3� Z|O�ᢇT��<^h����9\�#��N8�V�����AǷm�[sB��J@�"��Y�:�q�:d~u���t3��̪j��A
����(.�q��ѼjޱS"��bͽ�/cV_�Y���m���|���G�cYˆO�W�i��4M�+�il��0LH�z��z��JL����c�h�Q��ƗЎs���d��w���r�~�����P�2�Oq����o� �ٜ��\�\Wj��j�<8��HˋK�4�����eȒ��xt�����G��o���?v�c�����td3Ģw�b��j�*;����37��,�m�u�/I�&w��i�fLld����qԸ��T��&����sƤD�eD�v&2q���f`��ZsGKdY˲tMՆL#`a;�����D�$�@��`|�c0�C.�B�[-b?�n��uܙI���d�F��!C�������������p���cG�q+d��֑j	j"Q�F���j��Y�2��w��hNgB�>���ݍK����+�ަ�J��n?�88՜{O�w]�N�)o��u�s�����V�ݥ��O��6(`��F��`��D�!�_��s��s�*�k��hM� x��Ln�[l'����Ƣ�#�kM��x,���^N��`���qK	d�Y�
qZ�h�i��������d��%M���s�D�r�W�)��J�N�h }ѱ�z5� �=��o���n��Z)u���z����#�Q�ܨ�o<aVn��qKDܪ90ё��%[jx���'=�Xׅ���_�����U5�s�@z���!Y����5$���� s,R�.%�ᠯ�)��ѕ�;}��wMa����k���'
!����o=5��)���4���mlf��؞�>�z9�����}�y�Ë�[�!��I���Y�O������ŝE���W�ٔ�%[G��)Q2��X�A�E؛QD��N�[��!�x�#P$��U�if��u��ђ����Î^Uֹ�.e*{�Ӳ	� X�ז�b��R`���Mܪ���D���ϛw+����Wk��:���g,ժ/1f]���f,���zu���M�ԑI�G��Y��_�8ح�=d�*di~��3��y���
���م���Y�� �l{�O��|d�b?��ըIJ/.�{���*|6��F�^�6_OSL{>8��E�81ډ�bU����=����=9��V��&DG.g�9�n��v���|�����U�Ì�,�{�c@`��^,B��o	�!7�~� $�f�	�/Ŀ)'+��I�e^gBfR@D7���Z���*N")�_�F���� �TZ�[k8�&�:˝X\<��mc6�Dbޠ��7�ә�ݟ|��L�"�-�C ��h�|�믷���/)�Rap�L���8WPG0��"���ߩ,��:����O΃7��W4Y�ІiqWeнL�TE�����o�c2\��T]�Z��o��^��%@����
�M�t�?oXP]4U��܁�.���o\L�3�F����Jn�l�xf�����!��q��d����⣉�����2ѐs.�\�̆*�~�v���IDs�s�cKuI�y2�s�O���#�<�hGrI[���V|���,���#���Q�"{Zj�/��G��2��[]$W͠��9+�m�P�)	/��cDWsR:��b�!���n(O�_c� V�Z
�yH�eÞ'Zi��qM%�κ���u�(V���+�!ZK�����1n���6o���^!�ب�
���4�]j�<��uXZ$�}?>k�M&I|<�SR�N`5��K��7.�KY��OY�3�!�oUWw��!�������d����m��{���`��,�T�0��,�E��S�8ȃ���8}��eVqwdA���V>k�<v�ZV�9��q�"��.�˸�gЕ����������Ѳ�4��!q�
�[����d\��o���ҕ�a��-�W�ħ��爏����ӌ�Z��R���j��PW���
6�SB%p�u���{��%4DcA)�����0���1�a�S=ܼ��4|�ߗf*Ϲ:�H*wT��Tv!����>x����ʮ�{Oc�����_x�5�֔؜2����ܮ�*�JӃ��頠zW��_��`��h�Y���|����,yp�\�2:�?�P��r��R!����J� ~QԬz`&y�x���@�|��C�{�.�r���GS
F�iW�Pu/�fs��Hƣ>��^�M2�$�`5_W��&T����fpnȒ��PK��U2ꅥ�I����]���kn2���Q���Ht����fG}�&�J�!�?X b�˂xќ|�ׅ�Y���U\���2��n�<�$q�=�.bg���v[�:\�z$⣩&�-z��N�'^A7"A)����ؘ��$�����y+��u�{=^�FrS��y�OV�V¿z��g*��rtNx�ȩe/D>���Jx���հ4��0 c׋1i!�s0�����>�/p*ݯ�<�H���G!���UX����!��O}^Y�"Q��a��̆=�V� 
q������&���_�?g��P��t��<�N�? ���A�(�u�׈�Ɂ�A�:�ﯜ6'?��X�1Z_����E���<��oS4�n4b����l����	;*-�n���P�������G!��(ͨ���Y{�Ł=�$ʼ���q�-M��w�����ԇi��K�*��$g��.���~�9ԣ�I�bN!^.�/J�_ѫ��5���3b��^ƢC�1^�{?9yYF[*�ʸP�ϣb��)�
�#�.0����S����?��&m��|����\.GnӭB��EHI���O�];I�&�<b�M�I��'f�� �	wk���ڜ���5��֐��9k��b;���:i	SN� f)A$��k����D4���2 �c�F6��z�o�8�n�0!��d��¤a/����i+�s-���O�@�K"F!��c診���y���wX��Ji�,ˇ�FL�x�	uB���q٢r2�l��8ˑ����q�{��]p���[,���q却ۢ���`>�U�� �Z�W����nw�(�-"�n�^3j���c�St�+��~�m{�[�O�����%a��b;c�7GA�(ې��Ӝ�%��=F>���f�U��Q�jwd{)4}1o�%[��'��xv�T�N.��L5����bơ��M�w�"c���R������wK�%���Im�m||����5p�պZ������X�s��U��h���	�X�F�AHf$<�0o*��q�Ks��J�5{1V}�ݑ��rO0��%z~^�l��L�G�wWŸ��H���%�tE$OuOW�'�%Fl�,��ET�T�|����6�||��ۧ�z>�<8�U��?�G*�v'�(�� ��q1H4��������.��2��]�_���H�Q�z̷Yx�[4�df˶��-Hs�g�is�����׊�Y�}��❡.�䄼>�T�"Zq��.7�Z���CÝ�ho��%1g�~�zV���\���?wh�Ȳp�T%�Q_��ː���(x��#�k�S�E>ٕ��/�V�k���r�T��B�P�0�B���h;V�'aݏ�ǟ���wuOyC+A�?锰�s��`C��l#��^M�x��,(;��aU���P<��a�q���Ǜ{:FsM2�B����&&O�:%U��SU]�񅬻�B�ޒ5�At�ʄq&{rwe]~�L_�1���7��J\���6F�1<��I��PE�T+Ė�9�_��]*����;���qt�V^\�*����'��s`���HD�4�#$����o�����������������@Ώ֛�yz=�ͳ^���^ys�	��&� �n���E��5
Ӳ7�;S�W��Xhs��)Y2��^$r0�v��G}�-̈�Dp��[�d��ك���NlF_W<�:_�R{��b�L�n�"�i��v�ێ˖�gg�!����Z+�R�c��~��|Emˆ����s�A�)��ף���#u4�r���.�Ql+HO#{�۝L2�])ɏ�g��wl�.�ɢ�r.��:\�{y1��+vĜH���� �-��,�(��3n��U�M���'�ͺ*�'b�%��Qf	z��k��~U�Ѧn���]DLHY�I�%��Ֆ�B϶^|�yV��{�2� � O�=N���ؒ�:���ԙ܌�>|a�
o�T��5��_�D���L0�S{� !<�g�{��r����l����~�g���<\u;|�Tl<yM�&��1(��N�cu?Px��!�eS�����m+FE|�W�Ը9M�S�Wv����%}�v����ּ#�K(�2&Ȥ�ڌ�Y���lc6
�@��a�0f��W_.�Ua������)x>m}NH�.f�H	/��5�`n�ئLX�]�09�3Ǉ*�/¢e˞�"d7YD��4���2��wm��n�w�&A
[I4���K�˗g_�=���("!c{ĳ�s�o��~c�s���q�w����֩�#Emg�:K�&賆A��W�#�M�6��%�饻ǳ<W0]��1�N��"?c�&�t4��z5���蝥��y2Om��2]�c?,�,ǽ��+&Ed�x��f��״6��F㾆/ޞ!9�8xn餡GB)��	�y0�[�ѿ_��i�h���X\۔�!��7l�]k���c�����
�'��WxA���jV��ynUH'l���]���������$/w�t�걋?�(\�Gd��F-<�o���0%n	r��d����`���hc���p�Я�u�ٹ�O����7�t�rż'�j;{����x�@�h ����T�{�j2^��n��H�Ȁ?��;��G�[�	��ѷlZ�r��v�W=���,�нU��|	��W��)~�;�zj9�&�V�ڹ�	�Ɣ�M��2l���+�[#��+���7��iМY��.:��+a�fJ>��Y� �l���b�|�|CsssU4:�h�s�?�:�^������6O֥��h
{]��� �J]������k�=��r�!��WX�8C�*<e�(�k���b��{ZIB �Ȥ�'�{e�{2�������TL��5�6��A`n���5>�ҫ�n-%�倆&2�e2@E�L^(k^�Ѽ���(��EPM�
�_w�4���u.<����&�L� G�¹�:���3�!��cP�T�g���˘b�p��5�ՅQ�H�c�a�� Pe�F]H	�֬�n���HM�|�:1ԫ���MnHď��@-�Ң�K��a*�S�C�-�j�{��7�2�dq��X����ڵ����4V�`H��[yʺ�p��=��>M�E���-&C Λ������>tf���k��63��W�������M���[��1���� \�I�����A��E~%%��+�4�� *YW︍�n����� �>��UV8��������"���VȅҖ�2[ױ��M[]��e�� h\�.a2�K����$�c̀�^�R��*V�����i���[�LՖ�N���5V���z���'�e�z��GE�NRK�*J劜e1�s�� S5�U��OKd|V
�ō-v1:��,��ȸԘ�'^X�P���\�P��opcs&+q�q����D]KKhZ���b]��"w"��.�:À^fn�	YOXk�t����F����:���K�m{Tv���B��g�p����<�{�-���T�P1��rW��/ ��ܧ�g�G�
x�2����Z���"����mAL�(�S�㫆z��4+��D%�x��A�^�Z�h�IÕ:�_2�С&
�SB��F��I��(�F����YCv���?��$g��	�62W	�	t�l�b;>kr����4Xɰ��Gh1-���~8�3��!��i��ʘ98J���T��<4������Iu,�a���@��(�$+�Jn�ۊl�?��T���z�ZLsq(>�CI�Pe��e�H����8�����[v��T4I*/R�QrM*�ʹ�	��<���ڥ���h!�@��2
4x�]!�~��`�&�M�::���0�G�m4-�gOsf���e�����&����*��(�B}&Q9���9V�CU?�(fGKv�ƚ+s�Q���ʩ._t�9ێ9:X�9���4����tJ����Y-N���՚\'a}/Y�J��ժ<J�,N� �'=vl�$ko�c.:��5DS&����e��F����^�B�����Y�WG<]�I�:�Z$����8ʊ���|��I�\��ޝ���=�:ﺗ.f��t�!��b3(]���N}�җ,0��{�txM�C7mDݗ���LSAѕ�Lw�RT���i� ��^?Tj� U��@��t���8����俅G�+|ZqE���اS4���������6pB��&�78�4���y���[\�X*w*��a�+n�f�����n��e�P��^��_eцHK�NI��wo��T���l~q\nD�ݤ�Rc-Li��Q�pt!��^�Ǽv5|4�p�w"&�+"!���A_R��꫏�`'�4*���jų�+޲ւ��$���~�i���,I�����w�Q��w\����\+j��`?+�BK�<�\�yvLd�T��C��߷�1�T���qrQo:���ͪ '~�䗲�3�<~l��6.$o�[y���_�Y���|�n��M3�U�r��<uk?� ���B������VB=�C-cq�C�^�D�0OCH}J����~e�!��� �Z��s��ߝF	Q���f8�	�tG��μd Vm	$P�0��eC'\@6/�hF��{	�)�nVj��J���;G=�D�棖K�N�"�Oc�oT�K��K�h��FTXAESD��1X���2��;|�-����7Y k�b�'�D��*�Դ�-i./���gp�,����j{|�cZ���l�s�u��%�6�ٰ�,p/Z��LX��C�uH^9�6'�i���2}<�Kii!ro
�g)�k�N<��|�x�R2�`|^�~Vhs�Y/:�{�@�f.Z%�D}�i��nI���0L��|r�FX�>r�#cL��`Q�C��BWRv��W��0�u��BZ�I����jŷ)�أ���B�?K�xT
���f��
�>��jܒ��rl���P�uݢ����9��	]�Fg�^cR XY�7�:־-8}���+!xM n2����k--�a]ea{P}PfLd�J�Zܷuf?L<�Y����]O�L/�t�J}(p^^ �̤3r�Z���� 14;�`�m�3��p�ʑ�*ˈ�~��Bv�� �5�fFXK�Vsx�2�I���f^z��'V���7kV��>��
�{97}�7O{m�炘]���h����(�[;��	�nR�'���g\MF�� ���m�C����bc��M���`����/������F�'��.� �WFW�E��EAa}�&ݤ�L��I!pو�����u�)�d��ɢؚEN�il*=3�����83��˰��Ĝ	$F# o�YoV���×r�jdϦq�8ݸ �\ߑ|�uGq�;`[�v^�HMd������Մo�ߩ�Gc���̏]7����QFի�R�����P�!>��n��q�}\/ �t��`����1�&�O����|���n�V,dP���8��tp&���m�rRf�k�nҫeި#�m�	j0۰������o�mH���j��z��}MO7�7���������p0"A�Q��^�d=�њ�8���r��.�ϥ���yI���hT]ցǺ����y��U��^h.�r#ڪ�@�����B`���e'�ae�>1�7r�t�n��d �G�. ͹�X�l]ͲB�O
g�t�8�"��̰.�Q�4Z��@�	px7�=Ʉ�������并	;�rX����6O�ɛ��q���hn0���JІo&��{I9�}����T�3��� B���;^�gJL�H�肔�B�|9)���gfn1�PW)1��<d�y}#�K���ј׃&�'�)�!c�A�Mh�2 ��x��Ͽ�@�o��j�M@��X��2��qG�)��0��XP��z׾�6�[y޿EM�T"�I���lWlםtAU���6�1�R�,�O�3�]�"v���e��>��%��6�
p�Hg.��AVl�il����01~q^�NJk��lb�S���.���&��o�Q.��q������k��(g�@����O2'���� ���Hɭ�Ա���^�:�5ƿ�Ԩ��X��#�v{�<p�u�k�D��C*)�BuB���1T`(K�zD3��N�F-,X���.� ȧ�Z�ՠ��mǄ׬d(�`���R�"��Z���,���.����F�v���lּd��Q^,��$Q�'��aR1<��튙�3��^��3k-P���+����T��kǽ%�XÐ��䂆������(<��k�^XȪ�����0�jO�SS�ٓ��AúL{8�=�>8�7e����^�)���s�0/�׫�d<��lPV��w�Nbҏc�uZ���9Da��B{p�[t�d^�B3��H��ϫ|����m���c*�!��L2(��.�U�H��G�R΂�G�k�ёM�����Pu9G����������+�el��v���[aݯ���]�+�aT�=��yo�p��Dn�O�)������%2�� �4e6}o���6�=d�,���Ӛ���Fe[{o�4�/��>K]Oy$��T��8_}����E�W�s�A�`�5m6[�^�e>�u+�X3N�tfĔ��w�.!���}P��6��C���r0�-���Y�.[xH�?������K���}�6�{$���6BG�pw�̀m��n>����+N������]�\L�G�/%��w�|�p:p��.�Z�2�+��_�ޭV}��E����C��n�Z-Z�K�&�`��T粧U�f�9���3P���Naݎ.��nq:�5I�~W�Ҩ�3�4l 3k7N���n�\�yG����=���Q�xf���@,�v���0���0�},�q�jF�4z��b���<�4��	S��(ٔ�e}�m{��ǥ�(I	�D�,*�۩-����W�v�"�{(n� ��ߺ��vÖ�]s\ayo�'B���u��ȍ�f�S���Q
�V<�ҥ�ez�a*YR~��������(:�Y���$ɦ%�;�8��w�L�V'�D�V��-��C�r��Y�{xO"6�Ք�|���?X�<��z<ۈM5煥7_`d?�c���Tz|��i:0�۫����3%?���|0V�^[Z�&$˫l�?�A��?�RC�Ju��rt!�z�!�]5�z��	��s��]��+tn���� 1�>Р���އ�{n���U�[��w�-�;׵O3����^���X�;�N�w�_�o��ƭ�d7�O�n,Q-��&G%� �t��3�lu�ñ�
�h�a11)�wH��ʨ�Kŷ:]�Et�'���@�½�N�D�I]+��dZ��G|a$O�8���#��q#M"5��mX|-�f3�ӭOS�>��o-�Ek�2�f�U�%�Z�6���5ڑ�t�� ҩx	Pxƌo��|I�Ρ_%�hM�q��L����O���� -N�� ���8�cg9:�}=�8�/l{�]vM�N�6P�c�Zf���x�C�:2�JE���@?
'�}�e�eVZ�>��
sh�x��~����u-*��2��ƥԖ:��e/���Z�p�S���&���3�6?�ʹ�B��ٮi!�]��U"��m�픽���H: �7��R���k%j���m�Ff�{�i%H_nc��2߉�?ޮ3�tr�X�
��7�X�[�!?|�w*/� �ÓGwf�����󊵸I��I�n���fbDQ��j��ˢ�(�N.ʭ����V�CmCZ*O!k����=*&��I�w���
f`ϏZ��+�@�̈́;�b�y,;X��W�#�"i�'Id=z({�@���V�QؾY�:���XaEI����q�W�Zj�)P�*/�W��1X(�ɗ�,�$��\�^�ǫ����A'{�6!p���6�璃���f��a�H�7@%1X²��H1%�Hz"g>Ű���р�o�7�t�l{
��/����r,\���ɗ�1`3{�7�ӕ0�X$`�{�N#��|�����Z��T�@��*��)�FyY��<1쨪X�����,<9��Nj��ȹ���N��e!i�#h0���#g�P���V-`�H0 �s�rĥ�������^w�햃��U>����W>�;XrW�V8~������"A�i�A���{�^�У�*
��E��_i [J�ע���֣
��S��`�z{���@�2bQ�[r]۳s�0�)�~a��*7Ӫ���
���$�5���'DB88����s��7�� �Yl���Y�|���=�|JD����U��e!0�n��$�A���r 9 ���[\�>J�d��s ��.����'�::ؿYC}����j>}�{��pn��j[V!$��\㈎��em��堠v8Ϳ�� E������+DגּeZ�4���	O�k�f(��h.9���YN}�Υ_��3O
0��(B��ף�\3��T�y�.�w��|���Û�H,��5�l]Y�e�M)��T��\�7" h�/�m�*�׾
."���71��D�bu�HV����M�Mn�W��a� JvBTrQ���9�t6kD����[�uc����X��e^-�I���=�!<?�	 �*F�6t�/\./�b>T�ƌ%#�&���oSY�8�>�A���~�V!�g-�����6U'ɼWܯWC��є��|e��{�V�{1�NS�0T�8�,v^��6N��.�ŭ򃵁
��u>'����!���p�I� �~[��K�іb-�rNt��0k����x{�����^Ul��� �����]��&;�AW�\��!�W��9�`j�����C��0�m_%���>޼p�*{k$�V����v�?�t�/�cY�L��F?V�?��x�F�~Hȥ*v:e�*\�����s�j �;:�bC-� �H^��8Nks��`�X��X�]�_��3��s@��6T0מk��H�q2Ep�����Bf}�8�0�sͼ+�-L�Y3�L!����Gyo��ævmG�'J��oD��xQlz?I�+	:*��������	��M��?&��6��]�c�;)y�]?��C�����o����O�t^d�T�V�����E��2�֓�Z��żtI��"��v槹��j�.82I&XA>a>A>���@�1@d2=��tML�X��	\��  D	Z��)��?�>sY��V)���!��R���	�]\0���{R���5Q`�2��!G��׍@]�V���k����9�������B3v�I��\yY�������!u��Q�z��Ϻ�T�V���b��Yn��U��ڌ�.R���$��O�:O'�>�>N	�%ƌ��g��;�FJ?U�.��U�]�[Ɖ�i��F��5�R!�?%1;M�C��},�Or�ɋ�-BH[����
J�|(sٯ�Oe�Ҝ��G�9��(��)���Iӭ�Թ4/c�*}T�.�;��1�!�;��	��\�a<��늒���%�� O'���7�����P����Uy��"DQj�9�U�j��`�����A5�����V��,y*=*>����{���k�cQ��G�!����D�U8�M��ً���������W}���S=��S�w|��X�:k��yC�F(
�����="}~K�*��,cI�<d:��� �#���C�����c��7u��<	��qYu��jN��=������X�"��Y-_?�+�0=��Y��G�U#xH�n]�3`�YF���4\�^��؝{�,�
|��������y�K���**�J\y�Of��v�߱h��
��}�`����A��r5~�8�:���#�g���%}C^�
l.�����*nf�?�z��x���c�M#I"��Yǝ?P���S����x��2���+�J��E��!^*�C���x|�/]"���<lѮ
�!/r�v��9! ��DV 8d��njsR!�D�B����'O��(k��������hEf�����G��uxxX��Jih.�۩��jW�U_ڳP�w8�s����"��/)��ck$ +b��c���1�[U�1"�g0Z�:=g�>ĝ�����G�v3N�O�h���ޣ�_Ls���� ^$�[yK����yv֎_�����zerv޽1Rٗ[B����H�N_#�O� �x}��)�f���"�h-��k+��92�|:ܷ�y�i�б�<���\�J�g3�?~��%��F�7�Z���W��B����|{�R� o�NO����5���m"�x������x���!��Y���=*��N~^]~]�h�z-z[�~�՞�Z�6`m�-/CV�Z���̋Әl{����m�[5��� ���&�ن��F����:��X���%��c�QK������'W�Jr�[��sO��<����Vr!�c=t<h�jb�T��5��ׄţw���ۨ�Q���C��ړ�v�(��3�d>�����ю�S�R��9fUZ�b:AN���:R�)a|�]�q���	X�q[b&�[C���`,�T����(P3v7d�i}��K̢W���9N���R�b����a�N�,�+��}`���`�-����ϱ�1���4��2��ʽ�j3�N��80�mN��\+p�Ã�̎!} ���P�I�+˅C���Ȧ���hK�y1����� µ��W�fȞ�BAI��H�0��W��3�Ƀ�o�~m�@Ta�c�}���,��#���O�r�%�^�ro�П���{vm��w3�b��׵��n����'	�涴P�"F�,�D*ӄ�`�\�P�[K��46�9��]��'�#��hȭ X��^�=O���"��F�t��;�݌�.��q������܎R�{�zZ��ѧ��1�2v:E�w)*$d�d��`�ݡ�H���ifyYJL��QM̞��XR&�*<� cU9�)���z]������A`�J F_�C%���lPo:Y�P��9s��}�W�z@�����@�\�r�e�C���6�oq��"	FQ6�M�՚J�^a��=�<���P,x=�`��$�~���Mg��9D�'�$�����L�2��i�	��[t���cI�턄,	�I��?$�?��g/�1`�;����lЛ���W5���K娔h�ԟ֕PJ�qr=w�!#�e(i��0��v�[��U�O1�]�W�q�9�3n�wKuPn$���*����ί�%��&}���S��ȊR�:L�\z�S�*��"��g���,EۤG��KM{�\N�N�
��[*H<mNV }�8Ho�5�����=������o7y��˹�>���.�t���w�c�~#�mm���ѿ�e�Ɗ�{�9��&~Ɠ-U���e2��&j"H[G�`���`r�+��ϡxQ���h4��[�U�1/:1=��2�hֆ�d�ۺ����"+U�iUn��*2�R*5q֝� 7$�B�1p��w�q߀4~T^�BsZ�[���ң|��R�l��n�B<�C�
4)���[(��.����	ؠO�H�nn�4�?;P4g��)t��R	��:�1F��Sد�ÿ�=�,i�/t��'�޲Òb.��#2�3���'*��L��p�2/ܕ�%Wd��}�.⌞|�����p�RM�	�]P�<쟅��|,:�	�ҳߋ��*�8XH&\J�iX����Y�����(ޅ�iM<�6ha����W$S���>/7�C��6ʨ{��-v���������tp��<����b�(��Iۺ�SU;�Ϲ��z�����(U����W��24�RM(8����'���aȒ4^�m���n$;Bw��8�#���ɠ��_�GA4����(��%�L�\b;&�S���>W�"u:���Lv�`��T
����?�/g�u	j�/�=�����mX��>��q��$�}��(�pS)�X_*f^骖�f�z{HU�J� �-h��k�~���/k$�x��c9Ѹ�)�faf�
A���'P o�%��4�x��CCb��]���r�[Te�J�/Z�m��fm�1��{�h ��k�[�	�O��V��j�5���tt�>��:�Ģ��s!�"��y
Ċ�{�� ��c[0�0�>�h
�	!ǈ� ��0� T��χ��&�X���^}��=X�'[}c�lm��W4$�6�#��f�-����`�s�KK� nX���BM5�G���_^�¹���7���)�^����Q�l��>&_���3x�o�t�������[����[��N]z�K䏦Hk���M*I�}�T�'�8�G@����o�Z|�G���5gE�x�w8Xo�������W��y,"���P����	��<�R{�z+����oƜ�����
є������`5�����n������p�rݑ:(uا_jl�Ms�R�܀����C�R	e��!��Gl�y��Yfd�����AX�4���n�џ>�ʅ���pd��/Pxo�u&C	���0�>2���m�����/Z��H�&$fWz%����*�j�T^�}��d�_�+����fڀ�Z���G����Z���/�r�ܩ�#�M�d��g1X�>B��di0�'8�F�hJ��F_�d�H'�N[A�Α��.<�*a WM��⇙|�&u����\�@�2��f�����R�ޡ���F;�H 5���M��֤���M�E���ۗ�Q[`�vq��2���q�B�A�37���
P��G�Sj�b�1.��{;� �:�w@q|=w��ގ��ETv��i��8�*v����]x,��ZT1�s�k���*km�D�BmCd�5�A[���ȡ{�*�_,)�;��J��%��[ �V�ؒ;4A">X)�`��Ԥ^�w��������k%Kv��'��������:�$�A�:�}�m2{̉��TXm4����AA���0~r�ۏ��n �
�}w,�~���t�(Y4�)�Haȵ� О6�wܭ�Cn���� 4�z�T���C�ż�r._%�;��ǥ�� �j`<f��p��-y�������XlS'r꒓�dzx-gB������/lmR�Dxh�e���3���ߢh��6��r��gU[�\�ʖj$6�����+u���
:��R����i� �0!ڵ��V�S�F��(pmgn��]��;5�K%.�_6�-��$M�Rjp��!؇�Ы��CRo$B�R��]����_Tu{���#�5Or-)<�(mW- ��r���&H�|R�b�՟���om�;[�C��Fv�ٿ��dg�H�LH�0�͟��݉N��|ԉć�TK�a�~s���R4b,�m(`J���s���zG�k{�`�A�C�`���k�DE؈�T+j�e���-U�����P��|���l��W�n�*��1���0k�w���9�V���cT�x.CL��~�>%_�&�C�c��	��jΗum8U�@�c+2~��xn����kZ�XUi����~��Z�V�'��0��[�D1��U���m��lc�ס�8nD�(`
vp{���CO�l�ӳ��a>�ʜ�Oy=�1-k�۱"��LL��/�M���/|�o��Z4���ѬAԼ��7��J�>39�=����jR<c-�J�[��4��"M���b��{���ޙ�\7k�Ou��ɂ��]e�[�1G-3&�w�Ld����4�yA�e�bd �i�
��Z<�^���V6&dr|��ո{5!�li���5���-� �h��t�٩��Ut�2N���D��/���|��c����Q��P�~S��=���iq:H�n2�Q�	1���v)a�U������2�3���/z��Y�
Q���o���Ʉ�"�w�y�oDq��F&1�>���},kኛ`<NkT=��>.�ӵ�T�j�򱂦=�|&p��X�6�ag�6T����j\۵�l?;p���d޿*4��|C�;$g�%C�d����e�ySۺ�x=��<e!�o<*���Z���p��9g������t-��H�n���H$���&���Ɂ ����!�}�1�$��Z�_�E8��*�����r���:��N�|B£�[�M�:���}�X�Z ��R���K3����ڭD�K����@����� y�nD6����0�U櫰�b����c#�,�6�KxC[Z�R�sU�\��s�3V��ʊ�Y;�&;2�d���u�nմ��i�,q��"-����vba�y��s�$QO>��6֌�w�m�9�sn�x�b��r6n���t��[��AT��=3���w�߾�1Ҵ��sn� � m��-�0>�e���c�q�ئ�J�M���T�Z ��(�|�p�x��~"�n���?$��dgL!�y��ܝJ����4�2�DZK?�J�'j�-/�-=`-��vv��e�����u�>�?X0����2Ӊ@�T�N�|m�a��fs��C0�c��`�ç�A^�cg�|��2��bE��� �&�Q�cՐ�0�B��H(U�}ُ��Z�w�J��m2Jz��)��_ĿP�����p��/wd����A�0��p(W������WF��7��ȳ9+H�TV�� ��w=��]�D���	���Բ[��o@zV��D[���I	Tl����<%�1+�Y��v����=*�@�eK+��.� � VV��v�w�9>.���3���3�Oz�;�����/�"����Q��4!��ƀ^@�PZQ�EA.�&�zw%�%�(z<�Z�P�WX*=}_" ^�|;Ar���Ξ�{X	��U��_[��S��:
�(L��X6|�q�����nIdw���-\ŷzlpɁ�Ъ��k�1[J"!ϕ���`���+��-L~N�֣u�_.�ҡ&�e�o�����O�F��8f].+U�W���sʷ�U�f����GD�x�7̓D�����h��9�O�{	��+�"H`�a�2ڞܲ�IH���h{������:��4Z���^�B���!�y���%u�*�A��Xg��#��C��=����?��C#��p��������"�:0k���F����!R1�/ݾU}��*��*����� �\p!p�*�];�%����)KG����V�w��:
`Z**��N\V�x�"i�0��|��O�m�����ʛ�L�k����9�� ~l�ZU2�ˆ7��Œ-FN�*H�_�aL���2��P�A���7]��{+���p��8L6� �o5D{�!L�B���&�U!Ԁ���l�'3S)y~6q��x��������������hW:�K)��BLg��?��І��e#��ȋS���8�9���O��Z� �1o���8���j~���~6<1[�}@b��-�폸����������[Ԕ��Ӭ`��x�1����T��^l��ch*a*.���n�ڵ-jҐ % �g�0��L(�"���/<�,DY!��1V�v"4qA��	l���s�<n���'O���jd}��$���UG|z�+H5+��>�ȔRfd!�s�X�4V�Dx߯����vo�IK�hF�
]%���u����������en���Aq(g�8�a	�C&P{/�Y��7�M"�rJ [:RB��iժZ�s�O1�4�)u�)�����Ƞ�Z��3L��FY�Hg6��k����3��v&�4)P C�L�W]LB*��R��1�|�ut��I7�M	e
YRp�GԿē�5�½?����-7��CiX!۹�K!��%V&;h��M���t�$3���ƈ0#R��U����>�VAj�v��Е��Ǡx�9��˱@�S骍_�7-��`�VD@�4�gm{�Ü���E_K�)����謤��l�$���o/����>��!��YU��d��NY��f�p�A�'����Pp��I��Ѵ��{����H��?4R�k�i/��ZeqƵ�M��ʶo9mL��W��Z1���̞$��˃�EJ!2��g�;S`���Ń�����A��q�����_8[e��ĝǿ���+�����C'(@�4�ss5�m��ߊ<DU��d1*������X�˚���G�nm���Bf��b|c�A��ٟq�<7���A}9�_�O�ڕD�w���>�U\��͙D�V��j��BJu=���6)�*Dه"�l�'Aۇ�{gp#����� �	fY 6����J؝��g'���M�X���w+�Zd�4�f:�����Zt�����xQG�P ��/��+�H�,�c�q.IP0��&��KI��݆,p���}�Ks�O��v�h�Х-\��/ ~j3�k$�&#s��f�ò�v������\<ڲ:��������W�P���_��t��׺3�y��©]T]bAv�
����pc	����4а�ɳ舀��.4��r=4�^�AA�xS9�`#!�	{(�E8��C��'F��/yl�ęX�t9�Z*�[J�5�A��;�j8��W�u;�:+��O��e*�<������x����H���Ե����X�W�( �|��6�m��/�\۸�0��+6L�V܉��%�Na�T�C��%Ea�Y>�t�>1�I��B� �;0+5����z���X �3{�ɍ�1>�~�X�]�2��8Uxi|�\Ò���<�YsB��-8x����{S�IhC�TG��|��j��z�ƣ:/q�a���8W�M2'��F*)$�zbpl� ������L��>Or ɧY�jˏS	�0��rf��U�
b���8ˊ`	�"�i�9;�B%$ ��%�7HEIN4ꥦ���X�[\jnW�|�6�4dH+gg�^p'�i�� W�sQ����kB>����C��dE�Vm(\s6�0�*J�ʚ�����	z3h�6 خ�D\�c�hA��[(�3��K�8��^ �~3��2-��L�+�f�-02�OwtU���V �3��&1$�ڝ���[f'�U�*a&�\F���[���]��B����-�_�7bt~p�xD�Gچ�L��[^Tq��6��I��W��vS���Pk@����	.g�ȿ�D$z[��W��-(�$@��"�%�U�ܠ�#�j��j\;Dr�X�SAu��9��Y��
D�(W�y�����k�T,+����t�X~�Rŝ����|�	o��y�������p7zSnp��%�R"D�
���FS-��ҠS�Wǫ6w.���Z�~�� �����^I��%ǔC,_����[�ng�ȋLP#XF����<��;`9E���ĕ��<V�0un-�f�T�&O��q+���{�nQ^����B�y�r�K��V�*�EM�Y*���M��x�����h�H���rCz�!o;�C�j=x+֝ԋ��E��L�B�҆5��U�s�{T"	_/�A��0T���/�}=j��#��3��ͣu~���7AC�+z��ߴ�� H	y"���+�����"\dV5}�,������I�X�B��2�2j�bV�v�k9���)�:D[���߿^N	�u��#K	w���:f+�3S��������E���\vX�X��.��ȼ�!�[e^���4O�����KD�&V=4sJ��P;�Jwi�Ǐ��:�S�k�l�O�1C'Dlb�mcB�*���Z�>�:_����c
@ �<˞z̑�y?�:��}k���S	��;���SI��`&��$H��vd�K��,J��L�Zm��NWo:as��78�Y���Z[e��jb� ��Z��c}�(�g����Y#�Z��&q����!(F{2�<�٢=�"�R,��U�_�y�~}��5}�K��f�+g�k�A%����ƽb��A?j�nu��4��d��Ф�$�~y�H��`�⃾��k�������vJ�ksb�����H�}����r�@U�o{��<F�P��JU@`�|n�}Bْi�-�����Īs���-Ӗp�#��ޘ��[4~����0�jm;���CAߙP�'��2,O�'E�CcU�c��>h1x%�Z��������q�o�K_遶P�1�LZ���e4}��t�x��;-�."f�_��7�@�>n-���+�y��qr�u��]7���!?��\:��T���hFJ)�>S��o0����K�24=�������/����s��֫�ʱn��-�XT�J�{�#�w�~fS���Z� �6L6Twx�}�~��:�o���vf��}�ho��S����Ǘ�Z3�'ViuR�u�5��(n��/Z��ҹ�سf�y�ˠ�[�����m�����Y$�&���9<��mۘ��.zfDW���!'��f�H��j�zh����w��Y�VH���^����[������w.ۏ��~'�Q������(e��9?���ê$���É�q�h�;�F- 1g.���)Ƨ��Ǆ�XnVI�b�kW���7�y~��A:f������c�RN�^�-Q�	�ْ�T��H�~�`!ک�7@6�ȏ���Ȁ�Y���/y�����7�9�j�O�Pԙ�p��zL݊N���mB����kK�]�=9˅��c�_W��i�u����˂��>�K��,�6�5�G�J���G8/�Et�h77L�^���i+=#��?�E��)�ii�,�$&����S�OY����M�'I�ԓ�uX;:��q��|��9ܰ�k���0)�ŶY��5$����é�Dc/�	$x�e�/��MP�k�"C2T�̬��S>2���jH��";���_�Zy@.%u.���ۣ@T�ݟ\sGR��RHpɜ/�Y>�%"R��a���:Ө]St���[���K�u`���:g�VbC\0B�Al����4�'"Cر�������x	�g�w��_.����#���-�_��﬩������H:�/��W��cS��R�*�K�"�Cجeu1�D�	'�@K\37�d��,?\�eM�æh�qA� y#�����j����� �8�2_�����E2f@� ���)�z9�x�m�e��؜k=��Bʪ�n�+�P[�j4�ү����?�����!^	x��}?(Mm�h9E_���G����*5Ћ�>�& Y��l���/��'�0t��v��Wؿk�f2�� m5�=+�=	-f�b�p�m
["ޒQ����ʉ�R��3�:D���S)��]��W-�O��|WAhðp��h^ɠҸ�O%΃=>Y���܊���[NX苂Q\�1�Aed�u�F^��k�˕�i�.޹��ϥ�����d���}+��dOlF8M[^�0MC ���y��N�i��z���A@}��U�F�طѩZW�voB��9lW϶O�X�*eG��U�1���V��b��}.��zꬰ��yRK-;y��ڍ+V'���a���s7�Ě�?�|� �"��R��d#�K.�H�����'�^�`P���R��X� �Y�	��P
oB\�����j1�hߞ['~4�uo��5
4�>{���>���+H#���<�#2���v$���u�/�,��o�Fr=��)-��̛���k�����Lz���xxb�&��< �JX�p��Z �q*6�#������v 򅼈��T)�g�8X��yw�'�fl�V�.�?V�QZM���K��,� Ș2妆Au�q��21CC	A&E���.!��'J}����2M	t�+Q���]�b�}�ųHU�T�AN���{����#�e��uN��w��|E��l��D5bi�Yy�Kk������[�hOw�@&-��]8��ĳ��U�5Xg4�^Ӿ���$cMS�/��ԫ&�^��K],Fd���v��� UO\Ӱ�.�k�Qڠ��fp��KQ=j9��O����δ趸�Ǉ�6h�>�X�88$5�������O>�ޤ[��"��B!��x����T����	�5£���
gk+~J���͓��w�%��0�qĤ�R�#f�jަ���Q	����`�a�3S�i����^²��B��*�zB�5�VE����@�$�|fW�v��}3d�t��g�&���(����*5zF`w��,��ܝ�m�Ҍ���kj��F]��xP��2��k�A��9���X��X�a�(fCxRM�o�m�
7)������3Q���x��q& �y��3�ln ��$�C�c2>V?��&�{N;������$��%��a�j���P��pUr��f�hA%��k��ּ�olJ��68�}�Sm�"M���#��V�Q&�c�p p�T;��-�xٹE�܃�"Rlat�=����(�w�"ī{(���-���Y�n�`����M��y��b�f��k�����0h��r�զ����;	�z�����I>�5�٥��1�}��غ��YI�I�@��m#~r�ƌM��p=X����1h�@�ӪzR��[����i���(�D����� v>+�氭�9�=�C�b�"ݓ�s�7cE�V��q0�p��;4�iC���	�7�<H�iiX��C����'a���j�/�S `�/#&������K/�z ��|Mri(W���;8'@܎14(��VEF��3���^���/�W�w!�8B��g\���r��iq�fQ�3Up{�Q�U��Q~�f��A/{ZE�a_r�޼�~L�@�Gן���Z�:ՐK�j� ��;�l�Z�bP��m�6�cQ���L��z���6z����#��G���)RK�� d����jo��9,����Ӆ4��Wn�C��]j�T��v�o{^���F�^��R �/Hj�e�%�����3�~vY9�yB��Ft���^ѩJEHbF}�V_B��ո�%;�{eʭ�@���z�僵*Q�ƬwN��(#v�>�a�yb��L���i���/ b�t�F.H��r#O��q���_lq&|�P���SPzaB�3no��9����㇝�煛�)�?���B3���:<j��?��ɚ��3��h�X��ԥ�I�o��&v�q &�'6��8wwZ�87l�E�h@"<�i��zE>~R�B�4�������Lw��{��y��l���j͜���K0'��;\M8��6���E�bͱ�8�ˡL�+�0&�d3�R:���'H��Þ�^i�����GJ���& ��"7��D�=iD�_��/:�[M8�R�`��Z�md�@�k�� �i7@�^�w¢�����lu����5�9����WD�<�k���/���z��<?C�Kn�$���ޮQ��9�B�f7囚�HܝȔ��FZ<����,��(kއM��FW�Ǩ�p|c�o��s �*�-���of3��C��r�ltN�T �~�D��t:I�	��HӔ�2:��<]��"3*^���5a���1C��O�#$��?U��U�$�����LX�6���r˰�{V�h�t�}q`����� i}��)K�}+�qy����%�Mj3wC��hva�˖�jG0쁉D��_��/���Rv���4Dԣ}��?k���fx�G��S��szFʣ̓�c��H
��/���d��U���@Va�K#e���$�Ŭ��z��M���r���>oλ4!?σ�v�7:���(���=R+�G!΢�̀�A��f�
���h���F�UT\K����:x2���/_��m���/7=����{L�33;j��WGv�*���Q�q�˯��w��czo_��*$"�s ��+���m<
�^�@"��Q "�lz!*�@�[��P	H'.Q|�֋e沑:J�wۥG��S�z�� 0K�S���ac]�t�k�6�d��)�.3���#��r��i
P�h��w��C��_��N�y����u��W��m��N>����0�"3����ws����a�6�Xܳ�5�d�=��%׾���=�ow�C�,�ׅ�;�O���{z#�ܚJ��s���Z&]>�
�dZ���䲛���`�5	�L��*���2-���^��[ݑ·�n]������@��U}���JYa�_�[�:�*B��ş�����������(��'�챋������:��z=��
B۸@?���u�X�	f�ٵ�<�r����иà���޻K�z%B�<i�Tp)]��<Bg� �&��{�!@[8X�d�#����ryi��j��&u���5�m�{*OT�%�8M�w���dH�����n�	�x����]#7���Ka�Z��64��~3�2�l؍3�M-��O<to�ĉ�
x����L�1o_��˩1֗Q����w�8pc҈��3	��2�����_g�	X�j���Pl���<� ��=�k��	~�Pau�f�?��AmJ͙��m_f������#(R��������\��L@��]��X`��.�*`�Yyr�2�E��d1��XO��ў��^x�K�#>'�gdl�g��~�� {L�[8ű���� �̌"��_��gdu�U,��d�d歘r�uu��|���M�0[e�u&z =
�ZT�_M!;�+�X�e��捷��ғ@��g��5���fO�iJ��{o+Hv'�x��F���:y���	\n)��ec&���)�;%w5dp��A����:}nXN�?��?��?���W��ʭ-<�}RR��F�g�"y"�iҿ+t������<�m,�9foL�І;�<͂�ٮk�������e_�js���X9Ӯ���r�`���}�G�'$n����q�帐��?��Ց��"�����˖N��SI"^��ڊ	�����}�%e&��[o��,��'�TɄb��pr�{�n�S(�X|(V?B�2+X���})׶��K��/��r��^�屢����-!J�&¿]���]qv>��0Z"�ٔL�虲�`]5I�l�?�.�@B[*�*q�������P>�i�a�kP{@��Z��\7g�81�n�WC��{4�/�g�"{�N������U���pM=7�B/kq��h�������%!�>�3ad�,����v������р��EÞl}���6�� ���=@��f���@W�yؿ������$���Y�Z���a2��^�s����[P���������r�*٘B�LU��j�R J�L}|���o���."@�����G&`音�M=�7V�q(�w��_bl%Ɲ&���B�ia�9+�`�	�]����p�m�G�2�����<��fV.���"�1#��������8��ZB)y��i`O���J�l�[l���&M�4�UyZ�O!Q�Xk�R·�S ����y{V,���_�����%���	'NF��Pf����gI�������dd��$��$��1��4�w؟R�8�^ܝҰ���@8,��
�Q໘E)��TYM^7��dZŤ!����8��80��� 2�,�������zQ��!cWN�1{�=;k��W�F��B��0���� ����}zXY�����RĞ)}�ֹ(��0R�p���� �\�=����`h��!d��2���@� B��C_L[�C4���:��u���#��n;�c{��B��_���M���v�:��؁~;��rp3ݰ�q|<�	���V��8�mx�-:���u�ؾi��c�Q��n(�5�s@P�R0Nqs�4�)@S=�~u薉s3q|z�
��М��d�| Xz
��	��ӆ���~����=��#3�RD�D�"���lU�����7�	l*)����B@���~h}}�K��{Ժ�>�͵��O��X���E�lG�����ǀ!W���nOɀ'�ݪ>�	>ZǓc��c0Rz3K������2{\��L&�R��&����@ 6q@�^��)�e�*?�WH�9�J(+�W�i�X����u!?-�h���>K��݈+���~���T��/*����6�e��/H�6yr��Q؏�V��R͢�>��/�(��޳�X|��+��GZȗŠ���k�s�?-����ȿb��O�	���"ݷ��U8���7�um_K&7��k �H�~�e>`�������w6�Aϲl����cN@��"
qf}Q�����oU�%���o<1U��[""F�T��$>�� ��U���Bs�vX���Zeq@����"[_��� 1Q�%�.�����n5��JqO�׉��u�,%�O���Ϙ�D{Ati��v��E�����]~�����~5Z�������k9�%,�7�z�v�?���uzپ�����.v-^��싚S?�,
D(�ɰ��i߉Y%�=a�X�����}��o���K���R9VʪE��y��<��`Z��kz��mȥb��0� �Yq��G3�w���?������a�G9�.?ޔF�/	�W���9�7��1��A�z�G��0� *�-
 H�`�q� �+����H��n��L2�V�a���]�J�\���P�10�Dx{�ʕ�ߧ>.oo���8���m�cU��xt��5�c�d`���(��S-�\�ȢR$>���e��{�l@�cȧ���Ҵ?c�/�Ը�����L�[L�a�'H�P>�1��n�Fnh�gy���I_�:3+ �bN���IC���ԇM:Q��5�7&2ȃ�"��t�������9�g ��I��R�j� '�2A�ީ`�d'����!u�w��q�$?t�J]5o3=���j��@�hkHU�ps���rc����S�� E���U�J��b�y����6��Y���&Ku�#�t��cl�g�y�ؘ�n_F~ke�A�\;H}�w<�R����|�����>2�ݐMV���5nr��ԓX��d��T��a���yu�^�K/�3ſ���z`��h~j�M�����6q�7X1R�gIy��`�#�	x�MQ���B��G�a�lަ��/UɁ�";[�E�	��08���.'{�Q��f3�\v�΄5;�:��Q�nK��-��NN�s6�H0g?ex����	�H�j�?�np�ĩDK��oӜ�Z|^��G����9�ۙ��m�-J��i��}��P>�S�ū��A�-ĵ<��t��ΥȲ����x�M>�ιG7��C��L�H�MWa
�.�T �Mr��J�k�����j{�݇LrZ8|��F��� ?��h&Gh0������O)s�e4�l�Q�sS�0�YR�o^1��N�.Mll��f[�dG��8jS�$ǻ̭��)ʸ��<6rfg�`�E*���/������K�n>U��㼊�A�h�b-Ŧ�;�Z�4t���V�`���I�	ٌV:�r��%o�S��?�s�k����8�Gk�M� U4��ݒ&^�=UZ��{֋J��O	5�B���.4S_�Q7փ���G�D�o釨�����,�P�@�H�3���.j-	v`��"��� ��c
[�l8����;����ok���aL���4��(p�4����0ep2�)s[�$�k�>����0~�ƛ[�~��"]V�+os���'p���b��x&���jyH�>�����͠�Z�Q�
 Zg����F�(4D=�qy��!y�2=2|����K�����F
3y[��%c�
�2�$���v����.K���$��$������r�������m���\���U��9�����q�I-�Q���T/� r?r��<����W�"���H�7��; p%Gy�QU�`�J5'�����Am�=�QmfI��sC�uƔ?7k^�SF�D$:��^�_�ɯ��M�$�-�˒\=���]=��C�`I4!���"��콨)L�����yDJo�e,���b	��Y\l4/'W�a��ɠ��f��=<�0���>�{�IU�;�וjaWx/�ǅЃ����S)#�|�{l\6�1������=�Ҧ7������nX����7)BY�=�Q\�Ej�ݳ�*��{��[�p6Fm&I��-����eK$V�䘭��W�Nf�V���!S���thܯC���|�Q����|�oW��J�| ���F�tc�LF������P��i-aVXM��!n�X��d��]&lY_��c�I_�^�p�,pԣ�� (K�`�ʎ��y��x0�gR��M��ӷ��ՐI?��	Y��{Q�2�%M8k�M�$�,�5l<-�yZ�!-�/��-�4S8�Z�Ev
�`z.h|�5�f���6�o�D$�w��A-h���纅�T�X�ɿ���r�#� 4��]��q�#ŉ���%�=���S{���vd������+u��V�|��o�Y������$+m���Ƕ6��_��L7�(�}&ZY!�� B��&B5�(�:<)4�f�Ჱ�c}� ٕ��I��޳�3Ii���o���xD#A/���k����x�c�� �}d����@�R�c~��$ƝL������h�va��p>m����#�<\l�}�r��!C���]z��=/l��?��m�+[�����V�[]�@Қ�St��Ls��}�ᶚu�/�L	�wuỈ�^�:R�+�����On�OK��	�w�4�-�K�A�r��h�1��BlމF�����s��(�<t�����d���_��<)��!<�lS��"I�d��Pv� b����h��vn�<x�RƋf�)%I�Pȕ���d�'|�[%�4�������������-�1�9�ݍ/练1��qY7��XuQWH�ŷ�+Sՠ��r�BMh�����FW��3�M���C'Y�A'����(XG=����+������%_�񗤃���H�)O�k6{��*��~tQý�i��.�l���i&!����4q:��*�*����:��$
3\0�沏b����Ϙ�mU((,:�H"*x�v���q%��ǔ�._i�!2��>�[�ux�A�v��mXĥ���L�LL�ŉ��R&��j�{���kQ9�e��|��YB3R��-�FP �R>d����]�2��L2����1��o��&�B9D[9(�?���8��^-f���ҟ�L���Q�Ea�B�,�|'P���A��r=2�Epϫ��q[�]����k4U���:,t�ͯ�~��п�U���#qdJm<�M"P�>�f�Q�UvǶ%����?!� �_[�|7F�e{〇.Д�������PG{����Ѩ�ȭ�<�Լ��L|�_o,+�ت���'��!���5Y6���z{�w������N��-ܸL;UQ�H���"
It*����#�N
	�����Kȼ[�1�͆S*"Fw�jWVӔ�o:��@�l*��(��@Ǽ����d��T�7���J}�G~��̦�_R�+9�� F�*r�>�\��W?����,��an�k�I��J75�ٻ{M�l���c�����N�X����X��C��#|H�))3��}�	^��}�w�����r�6�w+ha/C�DO_Yc�i�o8NlJ�i��D�5��F�)i�}m���̴n{��Zh;]��II�9�����u&��.L�~{�Eܥ\���6}$I�����S��hw��6k�W��뗦ۂc�}K�AA� �>�m����������pPz1V���J��4�?��a9'��Ā��G�|��*z�G�!����]�n��Z�U��l��w��~GEs��e��o��e1
�E2]A�N��� r^���!��8�����~nZ7������S���c�'�WuC�9pHZoE���n=g����� g߿D6�A���P����,�F�[�5m\k[VS�e��Ш(p�qW/(W�	��$B�MG��4���O]���/hd�ΉέJU�s�oS�vms-j~)��r�Mf��|����z2��L�z�����]�&*���9�BIJJs���!LT��9:���������uk���$F3���FvD�u;Av�8�G��P��wqh�q��
¿����l^R��l`��<f{���IbȰ������ p,�P1���Qt�T�3Oz|?����(���+�X׫2y�ۏ9��٨�'YyC|k������a$�5k3�{ay��d���5�VK���������^D�����(�9u4�S�w�P���L-gI�[�Ͱ�u�K��Q/��B��� �S	@�)���U�7�91�a��߰帽D"�9�h�u9^$�̧/�߶�?�D�KOM�P�o5������!�}.�~S��E_&�SX[���]u:��\m2�u��{��{���o��k���y�Q�T�R�3�	@�B���"�X��� �����1�[�cʙ�b�r�ª��H{A���$��b
�_��-� <��u��c,*,���Chs#��Cy���~�#�C��-�4@�3�x�;�uם���s�ڝA���ǃ�����
cP�ڮ�D�}��Mz���W>Ȑ�˸A��v�Si�ѣ	�E)��	-s��N���(>k���\��:f�z��R��I�Bg���:3.c����۬���럡��3�o��!�RQ�{�*s2�ҷ
�5&[<jD���lU~�W�:/�՘G)o��Fl_&<S$Ӭ7����VƊ'���߿�	s�k�K}�0��9���/�����8*�A�]H�D�*6�,^��4oN����5�T���B�Cm�����$ہ��T;f1��o}�w`�>#�:�_�Dj�6(%�-@=M" $|H����&��+�����RRЙ��);��0ݽ_�����3�
�EI鼲�p;�jh�g���?LE�wǞ��˯"��@�.�~(|��?��G��Ż�H�9�D����a�,����Z�4rE�ˠ+�DJP�O�˗n�2y_z���+�����o�h��=�m��a*�ޥ?���f��A�J���I�b��]���� ��4�l� w��+ϐ���U1�z^s��N��֍İ���N ���������X(��+����@�v`���?Ye�z,}���R9?'_���u}"��%�ݿؔw��ΘN(N��+@�{�
	nE����ەT��~�H���ʎ�3�<#�ȳ؉	mS���܂��hp�S6h4?`k�DV�`�P����L�@������s�yna�a�|g?t��"���3�'.u�FǬlq�R?��P=6����`�cr"S��D-���n��`��c�x���@䙍7h؆&��S@үK}�C�n�=�%w֋^���K�^um����!�7_�<<��S��:|m�;�Y�y��^ �tu��4��4�E��s�#� ȇn{y%�Pk�17�X�H�SZmee�?%+T�]���2)�N�Kd�&D�{��/��-������H^�a�(�:lp%w&�ۤ���,��N������ ��s`�~��EJ�Ƞ]�}˱5P�q�
��1(����~Xh��AK�t�ck.-��غ1�}j
ǥP0�4�� s��%��-}W�R`"hTU�7`�Kn�%x&�$:��xgա�k�`'�&'���[���)�����~�W̯�ҾWd$�R����|������:�����h�����49�H���e.�7�j��RC�`u����f��Z���l�/�`+�b�稷ﷇi	=�m=0�g�N#�b���Y}`^ҁ�$S8(����� ����ja!��
A�w5DB\vW�����2Ӈ��	N��F��<��Vӡ��'�����;����|��7턮���c7�{��Sz�Y��L3��B��N�Tݴ��R>������v�Z�6X$ n�R����2�]�6i� �ü�7W&`����%��:fP����
���,�_�'Y&�a-%Y���o <����GlT��Վ{���b):D-^����C�^ls��$��"��/,�������`g�Q@�<ٴ���	#�f{(��2�o�K��5��9䞵R�v��u�,��EZ�8F*m���X����`N�GHu�
���*��0�_���D�<�u{?�!���������l���̷�����Dc'l������f�sߐ��7�'�Ϸ���j[hE,���~��"�4H�� Ld����?S��� �gӳ�$��c�s�+Y������z��N������nQ��-�GI�ڙ���>0+�'���s��"�Xk[���l��u�@p�3\�m���*L�S�Q�R�@(���FI:��?��̕����k/����88/ƷR���y��0�k^�o�_��zrqN/v���L[����y��b15Q7�܉��,�Yè�*eת���M���*���+�/�	��f��|K e�v�� ���}f_��@��;�7��)9����
���kEg�v��%�_�2 !����
��I5���I�����?Kݖ��$��%��V�(���j�(�W�>�|�=�Y���Rg+��r����#�;ŷ���f��e�a��G�;�����(��`�t��s�x����e�dP
ώ���(�D�@o�	v[�7S�Y����ڇ5hX����:LGG� �O	�^���CߢU������+O;���o��8nI��xFv�=������Fl���B��`:7�`�^��!}q4���:1	��]Y3��2�:�۹����(:�����XA��r�$����ο��ok�ήV�I��H���	��m���y�G��<��T�	�s\�Q�_u������Zw��,c�4H�����	5A�7+h����������g��M��.�w1�ҝ=?�l �*h���08������!�P�Q�&�V}t�����E�8��^�^�M����m{�\�m���+�i��N��0��`sr~�ſ2f�5���<p���� F��mq�7�3�t���5��+�O�/�d��]d�]N>/��U����p��W�;&������|C�>��"���xJ��=x��>���f9��hm��˰���NfD��,#W�jC�ɏ��&�V:�Ll�+D๐�r���gF���3���d���|��&k�{�_n�3G�ߛ�C��?I�I�m��qC�P�J��#�6��A�����l��0��0��*�X��,Ö����1|:���jw)����̞�4M����e����q���R��%5ͣ%俣 �'I�:��h}�ѷ*�Di�=���|�ۊcQ�����s;��R�ʚ����ML?�3��쟈��W�r���i�|��+�|�PB�(>�:�����v]�WP\t�v��Q�F�g�b������p){��n7OJbᏬ��B�U��{�3�0�Vxz���N~x�% P�/a�Oq?�e@���C�k8�oRj����<r?�E8h~�G����>^�bv�I/j�މ3+�Ş���,,�3��"�,}^�R�v���(�(�1�p���^�<vUw�b�v����c���B$)
����U��<���J=Ӡ�=����Gh*�AEyP�HΤ�.<�*�	8!0dB��a�+�lLh}�Y�B�zL��ڊБ���d�*�bNd����cYu��EJ����.hl0�%����n!bU��4�0w�Ȳ\���o�7#��Y����n=m ��R�O�^`<��Ͻ��fʛ)Ph--b�,�3�mN'ޯ:ݜQ�~ȇ���������6�����XbE	�O�BrzJt��Ks:x ��I�S�$d�}QӰ1�tթ�HW�x�S���M��­�U�-TN�G`����O��w�!ԡ��s���Ml�#,P�C�A\���X���h��7��G�������=�yE��U���m��mjV��v�V�b����N!�i����(�|���G��RbA�Wi��Ns_��e?8O�Ъu�� lþn���s,y&��'�VV��i@W��ˁ�D/���,���3o���36���d>����.b��Ie�a�4��~8JU"R�J��xT��¸I��t������Kŷ����v�I�?��hE�R��^�}&��]�m�����JrԘ�\$�e�u��U�]��� m%Q��u�a��E4� ���4=M��z�v0ff�S���{���^L�$�R%�.U"�����rAb��A�EY � �ܿ*/49N��2�B1|�&4��p�o��������b�>�ʰ�
�"H,���i�����R׻W�!,V�8�;���?/��lH�5��mˣnR��.J%�Yj#��%��O��P$(R�"/j��d⢷�#�|:<�����R���O(x-H�pyX
� �I�d3Y`�����Kz"��=m��&�ѱ7�*^�8�@��q�o�:9���<|!HvC�صZ�-�e�:�r]��g� *Q��"l\��@P���e�j	powV�J=�3x"�n!y(��]v�k	�PV텷-s���������Ӄ��bX���F�L,~�W*#���{��o�|��8�s�1����s��I�{�."��Zd�*��Rri��v"��5��͞SQ_^�����v�����!N@^��Z�H��𽮆�#��d�Z	)uД��3����o<������4Xא2փQ��g���N�W@�_�qFo0[�B��D�?�1&�RNߧ,9^ CG��2:.8 �z��MN����Ӷ�A�³��&��J��g�/o�=����6��y�O�l�1���Z$������,i/��"��'���I�M(!�l>3]�[��p���_ߜv��5ɆC�CB����c8��f�Qd�����	T�2��!�I�Z�N�-@kYNnw�(^�7���f���� gy��ڄ"rZ�$^��P��� ���	��>J�dm��D.u��ϰ������{Gl1��CS�F�g�5��[���5y�]e9��V���=˵�֤�yr���p;�f;�w.� �á�4��D&_[�@{;=���"�ӈma�"gG�=�`�=0�B��*hJi����X���I�]�TP�Ep!�����12�H=�@ƞ-�f�6�
`�ZZ[�L��Ɂ�K�\j�H!HÂ�ڤ�П��)�%s�)Y��k�,�P^�"�E��%ٯ��x-!Kl]c*�-�grk��1���R�\���KS���[�.�2�m9��+��Q�I��=&��凞9��~�w����S��������5�<����d��y'g[��]$C��g�H�j��Ն�'������`���HO�3h�zL�*��g�-KRv���o8���T�j7^�LѬ���rw���̠�(��{�%k��Ϥ�`��櫟���IK�?-k��۔��0`��B�uHj��v�w;>A�W�v��wR�Z�vc9	�o�ӡła�G��НGd]Ye	!���b�>'x�m�ۮ�p�ze�?R3�:����#�Y=�I���4��	/O�0�����O�z3�ݪ`�*��>� ԊJ�稸�;�w�����eǑ*��7�e���r�� �\��ن	��oSC��,��oB�{^ap��^�H#^l���2ʍ���D.[|P�j�,mL��p����7��9�WN���6P�
�[m���̯佥$�+\���a4!n�����Fכuw%5�%�p����m�Lxgu���&�ۇ4���S5�K�_/�k��i	�o�t�*�#Bq�����-�w�E
%D͘Ğ�1wQ!~c9�ֺ��)VĐ4&����q����v��ELȕ�hc(F�`�:���)H,���⸥l����Ʊ�,�W9�{��O�e>��C�q��Q$
X�ۊg���Ւ�ڶ��O���}�5��tr�,Zp�nS��"��m\ufj:<�r�`���9�F�umz����1J2=�(֯?�K���	4L�9,O�� ��)w��o�ҝ��ȱ2��f>�U�B� |!b�z*9f��FE0N�x�VyiE�͚U�v��<|��\[!qV&� ���ᰎ{�<*��h9��ҴvB�����g�bo��WІ����]��A�c�))���)N흊��	@�8+(�B�j�}\�y���6q.c��M�ѵD�;Y�T��\�v�~�y�r���>�C��:cm�ʊ�����l(v<ߖ�k�v�ނ6G��S�R�.��և�j��iF�5������jST^�(��P
�~��>�}��
 �f�8�����"�q���Vǽ�tm�dx[���#�PJ8�&�ҳ�pU�t �鴧^���$�炝-'�̣�v�/W/ᨾ����є�,��b��c
���q*��YW�f��O�G��� �a���J�	���̄F!���ˉ�h�T���}�|Fw��o#�= ����]��n��иelԪ� \��I�5�\�#L��Ñ>L����3��m��X��̴0�V�)�򐤧Y�s�8u��>��d��}�6�] �����j0>�|�VZ��?{�����1PNOC���C,�M���%���������=|')7|_ ��J���;���~\�}f>������r
��m�p{�$	�{n��K�e�x0D��+�'�wF�G5㎊�ݽ9kyj����_q#�D9�,V?_�u�o�*��G1��<��
-�ieY�ֆ��ZZ����A�������lL	�����c�XQ#��<�g��0�jN��fm�r!��4�9�Fs$D>���%���4gA�iw��t5Ɖ���=߼�Yht�@M����y��e}��uy;�%&��q�*r��$Yd��HG�?Xϓ\6 ȉ�CI���n�u���1|C;�Ud�z���P�ka���Ԓ
5�;L.���nV=���"�e�H��d��y��/}��kN��x��b�fB��|��Oda��h��K#�Jɒ�fRLW�-i�TF3�c|U�����#��C�^8��J�0�������%��ax)�����������N�&qAT~}��1��*��X�N�K�͑Z���<����_�
��m�$��9E(��"�0�G�ǧ;��ZW��X-(�j���޹x%z�ZV&4c�{��C`X�/�vR�2���*%��N��켞j���}�_�WO���xAU����3&rF��M��#ܟ��>ځ�ӫ<��Tt��i�)����*,Wlbw[`���+o����{��'�T�"X�f�zM�SZ`�b�̧I�<�)���aϑ)�"��}'P��s|C�6�n74�e\1�ʑ�%��*C'U��	F]���lw�O#��=�]2�x>g�C���i���>�u�y�d��O&�Ԑ��uV��P�c�$f�L�Y��X7i>��I//I�m9#%� �T��c�&E�7��-���Ђi�_������S��S���0�tsC�a��5��=��(ǘ��� ��6UB��h�±-���F���$+���.Q�̻P�H�C��h/�f7�׏0��;�!�f���^�{���m+�g��𤗂��z�F�w��W�W�S4x�bA	�L��.w�7�vK�7/{8�@��d:�/~��	Y
[�X?I�<G���S��=�C0J?pI�a�M��#g
��-�E�58��o��ZE �C�
j�vHK�_��f@5��z�Cu���6x�,[���k�&�1J-��̾w�g&�ߨ���h�I�����K�dE�5>�.�u�����r&���j��Â�	X�Wt�`�D�4�����HJ � �L�Pr�L�)y���rb���p)��R�	j<��$�S��M���,�~�6j\@�,*�f_�a����5�Q!:��\�
Й��$�TA�-�<�䰨��2	а�%��;^"�5Sr��8��W�G/i��7�'����B��Td�����$�n:���Mé×"L��+�:�]yw�G�O���Ho�PMS��.��1���H�8w����?�h�}��_�u��m�	�\�4nK�cΠ-������7F=#��wi���L�1�#;-߱;�u� #�i�$�h�(�uc���Y�&��.F�N��>�=U0�49� ���:b�}�!��꿎�`zE�m̌0bɗg��F�P�gh�,�A�TK+�b3����Ƨ�*'Y/����§q����G,���@B�S���Z�VA��#�4;�S���EQ�Zt�F��a.���5P���ڼ�{a�=�鸃�c���y��C�`g5&R�8�V�cD4�!o;�;�S�Z�NLa�=rpk�;�dj���j֑��{3��9�>-֊���LƳ��q��C��/d�l�*�������|����!�����0|x�1�3���}t�I×��$u��1�]FC�`�g$��,$�vT��c�+�Ù7���&b��2i��H-���D����Ȋ��b7x��j�:�[T�95כ�l�e=����TӐG�#�Z"ͺ��׾H���Չ��;�l�N�_�W&x5~���L�N2�<�̎�woТ«aw��i,��x�CUxJQ�fW3��S,��K(*�Q�7F(`\�ඹ�#ET����/GL��F^�g8�9��>�ٵ*�ۄ�[cU��ONϻ*i�'�m���cH����6��x��%�tT�本��2��t���>+A�����e�}$�
/(v��ctf�X������tc�ȼ)�x�m������=/��l��KQj�j�0��W�M�b��k3ݑ����"�\XɁA��}9S2ߝ���	$�V˯9E�p��K��2�l��E�pI�yE��	�l�Y�&=��s��4t�cc)jLqA��V{"��d��IU"�Z؀ޘ�d�&��6����/������LC$���!�y?c��L��T``�E�vO ���zT�X�n]~�2k�kB��ش��	����f0ۭ6�p7�xE1���������w'JӀ�I͝?w��'z�2�HJ���uk�;�
��e���R&G��}�ے��/m�<]�w%R���i:{�#|�R�J��U���Ţ)�$����V1��'��}��ńDCh�''�'�����T�2��U����g�)bZ�~&~"����������qJ�b�1�ˢ�(��{�x}?��S��;�:�g,[U�	!o�S���OF��3fT�:!R�a�0қ���5!����l+|ΛS7���Kg��S5�V7o�{pX5�y�phQ	Z���=�S�����l���9rS���dhE��n�Y�X[�o��[�+�p��\.����P/'z%��C���g�oXꦿ�xl���������u�������8���}�̨� �П�궧��A}�����T��qo��so�����c�G-�dT����C����^E>f�(�0�X��!"Â@�1*s&�;]��Xk�I�Sù��:�ʸ����Z����n>���,�����.��V��;�`O�e���{�΁�Q!��UW�c(�=��~Mc;���P��G���|�!r_���I�b��x3��3,�F]�ǌ�>�@օ�e�u��q��JF�M ��-���gg��ˆ��ʆ%X[������ �M3��[}��;�}QCT_`)�@r'O]��� ��?v�cV&O�Oc��T��p�W�U[�_>�x��Of"�+җ���u�Oɛ�h�q�����J��'�Nr�̺[��dUIq8���=�;ޒ+�x�?u�v(�틔?���s5�`�-���2X�1y�N��0�a�}a׼&� Q�{QP�?�o�
U�#�E]V�[�H6i4�����7�ۿ#�9dc�6��[�i[�0Я�Gb�G����X�qЁ��R	��Y��'�ɺ��V�au`������ϕF#H];.��)�2�a�h�ν^��t:`��ck�����~<!�0��r��]��G��t ��dq��q�Y&µ
��N�+X�Zo1������Vq�Ut�A��p�?ϱ���X��,��/ �x��۝ۋUrJ���.e��ߘ��;�=�)O������߳ݸb���ݤěI�9 �B:��\=�L�Y��V�?߰�r�!��<��!�m�O[��t� "$F#7V���� o7t`U�s���N���a{��:�ޮn� ���e�M%L*%�����u�ۤ9~�*�;��$�|���n���6��?�<'z4c�����lr�(?Q�Ĉ�w7��bn	ԤWᇡ(*���e0�#�ױw�{��y��;�k9X5z��ԯ�N�ظ��ix>�w�/�^�s��D�G5m��|���@�-{�|��i	7�fZW�P~4�.JR���uF�Q���H���^�o�4ͦmN��-�l��R�_���ܘOJ��?��uN�]8f�'�N�=*��l �<]��48��o�=��||,W��;*�-��`� �%�6��(cP�w����l�x�$B�g��ԭ�%'���3%�L�1�^��J��t_XY��1!	�J�O�:{a�m���6�N E]�n�_�	I��G.$k9�Ktݠ�Uu�w�H�q�n���%��V!D��B³k����*����J$H�"?Ֆt��Mt@+]s��C.��{y1��޺m҃�G0܅ O`��$̦C�X���Ġ�%����`r"���5����-Io��| �m��u����"���Y��v������RB��D�j��`�H�hkO�����tg7yG|�Q�ꐽ��x�ۯ��_^_�hu��z0SG�͙��yN�wR��G+���9����J-���]�sx^!}�o���k�	Mw�iڲ
�\��͐��	P�k�.M�.\�'N��鋹��h���G~�̓��մ�0:�dWS#�AZ�g�fʿ�pw1��Y����3�b�<��<��u,���@,h��7���8���
^I�����C<T��f�ar�����O�����\�pyDN�>]������46��ȝ�io�4��-�qpV�����z�H�&��*<1�1�^jC��7���~��~���n
��+��ڛd�.����D��c�y2�:����rѢ�� �.z���25�qd�K>����������v�^o"�ͪ|)g��2Ts)E5�Q:=����yx@L:�d��u��A���w���ѹQ�fZ5�Iyitp��xf/߉�0�}9U�|�=���q�S~�/HD���ub�jPV�X�ƄV)�Nm�cc먘f⪋�p_�����谧�`�!*�5kz0�i�	uō�P
'�;�Vp��n�v�@�4K�3Ӏjk�~I-)�Ɛ�8��Jnс�_�a�#h{�髮>����Q��H"�YX<�o�p�M�ƾ�'|H�
|r�Q|��H����e'�xw}�=�)�t|#[��H�U���\IOr���]G�FDKף(�Mɮu��+����5J~�CFK��Q�4	�K��Y�Ebc���n䏭�r��+#�P�d1���r�cq���q'�e�ձ��[Ց"!	��F��P��&�����?���=nڻu�-��\zU�eGQ������F���u���w�y�
�-�Q,� ���U����( ߹�V��*�:F �V���O|ޑ=�:�%%���u�d��h��D��N�x�?!4'
�Ѭ�#:&P�fF�u"�S��������lv�C�ce�;�n���L�~M������ {�1�TI�#�+��b�þ�$V�2P+]SS[��0I}IR��d���!�R���\�}Gp�
Ћ������i�~Z�����W��������79kƾ�v�L8!fh��;��u�5M��25�Ҽ�o��p�OkC�~�p�!�G��y��p�EӨ�\i)Mۍ�DL�XFVk��KS Ò��]��9�ye�
_qL�YPW�@c�Es���.��a���4����}�f Έ������V,��R#2�)y��2����(����#>���K=����5��$!�"��f�m�rUOj:��$���.�'V��I������Nc��t�v��+�����F�!z@ 0*F?�8�(:zt��r�[�qj����G���7���Xe��x-ЍT��)�����%5Z+%�tT*G���h�h���|�7����Q����?��dwߚ$���K�a�|(�qU=Pb0=K�6h*���G~9��蔞@�/ǔ��ޜ���d	qFcUT
���elE�{Ȇ�k�
�.�\);/���K:�HUK&7[rlȝ�����Ӂ�=y�`�˦j+���9������ux?	
�7`Je��*��ՃQ�G����\����s9�� �%k�w�5��6u�¼s+�P�)�Z��?h�3w~��3�j�8����+��O�.�����\�W	�ܮ��N�r-m��C�;������Ȉ�����E6�x���q��i���2�d߸|D>��E�9y�#}E�В������T�����cm��Ə|8���eJJܶ���n9(dͷ?ӿ����vc�m�~yb���9^�+��8t���W�"�����-;⋌����N��?�e�ɒG�+�EHǠK=UQ��t ��|�R�~��>hO'�>	�J��<���"� �}O�����=�Q�'E�P��T&�[_�	�]���Tw�>������	
?�+�k\��]�O�_��۞���� g��Ԫ���*��mL�	��ͫe��Zk�<bAD_�"�g̠��(Enf���b���=�*�PRZS����d< �[�Y����C��D7�*���y2=���D�T�i;Vn����݌�܁�����n�3���[��6M��<�ŋ�>�!�o�J�A'%S+g���c�6��F���FM������Ӓ�=�Dt�-�Dy.��`�e�k���	_�5�9���K��9���*������(P��:'w�t�%�w��"֦���t�|�h� �G���J�؆���.q딿�o�c�]]ۑ�|�ٛ�n�h��`�fʝs)���u��-�on��m�1����
ϰ>\��3����H	 E1�l�L�j-P��rT	ZeD�=:_�f"�?ҫu"N�J�����6J���҅�:������X4�8�0`T���$[V�Ҋ}��<�D���Td��C��%ǭ �#�� &r��G�c��qM1U=ɡy|\��BGc_<�	����N;W�T�s�a����/���z&q+k� \���RF�d��+��{��e�0$H�MG���p&����`�	_��bª����D<[�_���-�)�����F$��c����+��+�G�P2���f�U"a��������\�y�ǈY�b��uNѤ���%�圽x̿�B����gÏD{|I%�NG��I�X5�eS{e�E�r�OZ�
ݕ���Ȗ䣎`�>#�Dř���x��9��}-�w%q�jtw9t���t]��8{��t��Y}F@���F��pr�l���6���<�U[����*��K�g�Y,�������N�Ğ��5gh$䈰���ö#���$��.÷�!���{����\��p\Q۷	�!�.+_�c��*Af���_"鲴�����8�nv��#؇�"�HoWܥ�x�Z���+RR��HL���ln�Gp�;+�ĥ-��A�Je}�����9��S�O~C0�/�;�L��V���=�8{�!:�:��r�{�|�����\��F��Z��+5�4������2c�}�� zX��mh���(sʢ�T/1��p�Ȳ����!���Zhf}��uC�Uܝ��rB
��(���R��OY�V��1�=�R2V���?V�����~#m����$pɀ�Z4?����sH�Od��O~Ì�;�Eab������IT�+�������ɣj�zO�&�U4�m�ՌfYأ;�҂E�"���>'B`a�U�%/\V�?}O;����C�!X�������I	��"r��p<e���Z�@%#��O������g���7̅j?��r�Ơj@���o�q��<3n[�� m?N���P��6���y<��JzQ����G���R'��� )́�����ɳJ���~|�m^���<d���^�ȉݢLk����ӵ�_ՒI6[4��f��J�ģ(�i&�t("��`�-�t�����3���|��A�y�YG�[�r�4S���(H������!
�,��� �-4،<jG�n�B�G e$4���0% m�|Z�WF+���v�\�\�B�;J1�Z��	�=�¯�b�H�v�u�y�����;+#(ey��&��:m������U���=�� U���E�=���-R���_]�@	L�f�o�,�p(�ߎ��M4cojڱ`�ϠKD��PIx&I�l�e{�_*6|��0N,?ο\E�V��g]��6�����(�v�7�Xk��Vޔp��#���` ��d�����:3�afQ n��wΗur'u�Fڋ�-��E�:4�ɷ��ٰk���^��!�-\�h�XŅ���:78!��b�Izu���S)��k�8�?-F�p�Y�{cFq 3iw���҄ Ԕ��o�A{��O�D���TF�jg1�LJI_����&�����˯5�"2����[�kD~�{K$͓�����i�ē&�ܡo�=S�`�����g�W���QQ���RحHr8s1�9�O�,�;�W�u�m�o$n�Ж����>�9��Y�݆�J2>�V�_�Je��G�tT��YԾ�D�����{��mZr�<?%��r���� F��@;�c�\r���v����@�¯��M�q�� ����*p�g��HBK�/�Eիr�d|���0��-E<[����f2���F�Ž�ۖ�׎$��A�j�%���<�&� �Ys��L1sjS�����X��ǰ'
�����*ׂ=h��C���Ď�yc�sp�Zpz�� �e ���ؘ#�w*����=��ѐJ2b�0��f�H�fİAS����i1OQ޹�c�a�!EBNO��Ԛ�!b?��a4}YZ�3�
�uc�EN�j�Fݠt����	�+���:Ǫ:��gܩR���ozSO��iB=>+y	C�L���Ax�s����H���@g�$�(Ҋ�/]���z���כ|�h*�1�	ȉL��=�v�X���cX�_�h^1G�lM�mh�O�C9N�u�$=����	a�C?�͘M��w�X��G=���w؟��y���\p�,��>�ň"a`mm9J�$o�a\�"J�����M���S���#�����W�
��ͤen�Hх
��n�K�< ��F��)t�N\yU�e�A�T��V���"�;�-�[���9��zu�G�9�[{�%ci��}`�꽬����<e(��G/�����b��ϝ^�+N���m��!C���$� 0��G3�|�P�gH�1k����aej����n&H����F����=��n���M$e����'��o�_��������(K���@�(�q��a�;W.�C��m���
�Ul��V��SZw���ួ����	I��i�L��^�L:�ʀ�S$����	��n�<�uV�5RN/�2�k ⑐T`$0bJE�#^>I�ʫ2��+$�q��+�=�J`���i�ӝ��[��;�rRU�,���ȧ�J���O<�8ǃ�Y�ߜ ��X�R�4��^�RA��B?��k*��J|gf��]

n�F�Je��uD�\}����iD}��bcz{)Y�Ea��L%�,L~͍-[@ #��PF��64[C �I/2D޲�0l���2�dH7��~5��&�M�����9�5������\��Km�� ��	�i� %	�����TT���ٙQ< ��B�k��v
3���*{H�8�Hb�41�������\y�2������ת�1���[����*ιn9^�x�����՗�!!ZE
;�;.��4���!Ŀݱ�g�6���в��BuYX���vμJ���&����8c���pi�����/`�DR������R0�*0��C˜�aYbU����)�Ɔ��I�H�vW���Ӆ̡�z���ܰ0qcF�dY�%�έ�We	�:�� [��nEݚ��� �m:ǈ��u���	�(�f2z*uP1��2f���=��ʜ�a�[��T�N�0E|�ۚ��$=�貍#�ܞ��[�W�hV+��34�/�ꜩ���~�p�m�u�4���S	%���c��3�7��5G}o���%"u9v�e�D� ����	%G���5���á [�"�Ώ���#lZ��j0`+�?nJ�w~A�<6|F)嫳��g� C�Ư�6ƆOS��� Eo�
�|�W������&G��i�(\M����U��ѓ̜ ������etb`�1K�By��=�7�%�L�^6뮡� ���,dKW�s��O��RZA4������f�4͒��6r��#���b�np�n���үG�X��4���E-�Hb�)���G�nedb�x�h��Ɇ���uB����7#��_�l��ݧ�n��<��%j��JQq�K�|8�ԕ<�`��BU�[��ĥk_��i(����(�Z�Vy��)�Y@���m��6%��$� 2S��غ%�d������v���Z.�u��$<f��~�Z[��i�L��kO���(�̼�p�\7����mm��b���)��l�!�Z�-�ل�!��sB�gCW��Gs��]�[�>@�.m����f�7��֟\��F:�ʩs���<��rE��2�%'[�+&�Q�N`0SE!�E��+�'�A�N����t:XV����؜�R�hm����q�5dH���!Gr����'���|f���y+�$WB=�
��n6r���S^�e<���B��)�7�ʯεb9�ٝ��ǣj[-�]S'_�[��w����b� Z�����!�9��C�{Z��Y֘���H��b$������G�uA�2z ���mo%�31�Y�о�������O`�R2���$��Wiw<�U�����S����Da3RE	�=!�4y����-�.7��m��|�P�\X*M����Kb&d.u%��!�I�c�A�3�3�*�����e"�U(2s���L�`bEP�0�)2�)�o�#8�A|�u��;4���h��6&��=��8<���A�ѽH�e�>�N�!�䩑obS|S�����1��.���wʶ��i'�>J΄�����������ej3}I���z�
T���[���^{���%���&Q����F���'�R�n7}�O�u�+WV���SOn��@QUs�w5��#�>ecBdE^I�(;���tGu��S���_��A�����$�wk��k��h�Y��1٧�B)~��~u{��~P�ݽ�q��$+��e�T��Q��ʬ�v�x]�MQS+�Q�,�
=iuk�1��Y <j�2��P���7��r�c;�}*8�6���� 檣�E-�}J�qh,�"7����G�B�f���I59�Y>E����$ؓ��a�<�p���_i��x\j���q���N�σ��KC(�< �Ч�����>G�Y��W��~�l��+�<N��~��auy`A�.59$�N��_��7�jË�~HLm�i#ΆΏǚy�L׺�[��<�U!�ɈޙP��q���8�~�b����:�;}����b�t�l@%��I%/�����N���4cm��}�uzMi�F�v������ǎ�m�{�����y���W��{�w�]V��j�ܴ�|!]'���-+l�>B�xr�u��CG�r��1N�.�	kBT�B`6��A�B��l\��s��#����2+���i�P�Gd�(��'���t[�lp�6E�Ű�,(���zk�P�Ǳ?�	mb�u�`��i.��-X��1%:����9J�^w�I��	:L� ��͹N��Qڏ♡f�z��)��t�N��E�Sg�@�-S�`	�C�0����>���y6u�`�簤y[C7�o7/=;p�z����C��&��;�E�?��r�]�yK����6��r���,�QfJg��Ck������#3���E�X(�)eH���6J��;��Z�f�	�O��D��t� �*�|"ہ�[ˡ���b�J��=B^�,r ���׏mެ�&�T�	�08�P>抺 �{$��#X�=?@o������r/��)\e~7#����EZ~��F�)����(�-�}�����,�*ieU[�8��HWR�5�J��oP(�M���։ӈ��I�A<5s��)�rR�.`�L��xAz��#�?2T����6�^M�"$��pq����B�-�8�.�-�w�`�T����Z�v��-=sUl�����������@,�3C:��Q��Q��$�+褓[���7ݥZm�c��X"*�)��Q���֣��4?��_�V_�[���n�E�@��L��F�D �lQ{��e�=�����r��i�pit�vk�^��@�y�bS�lB���ܵ��ﲻ�o,�!�͂L���(=��T��6�樲�\�tV�����Ĝ���(�1���/�(`}� |��-���|c�r�q�����t��������Π n����%�B�	'� 8��{�1��9/���x� ���]�8t������y;��,�N4�zk�'fK�Ԩճ$S�ڕs���*?�9���!�J��٤O�Fv�N)��M�<N-s�Pƿ�V~��$F�6�$w�F��|(F����g'=颏4����j;����P�ﲼW(U�A�1-���z���@�˜���m�I��Zda3u��hQb5y���O���ġ����ajޤmbj�����v���{�Վ�O�y\?�Dy; �p��-�1�Es|c��K��٧���N�u�G�w�j:��|F��dˁ賈l��Us��0�S�'0�U;α?f�������w�����i��?��hǿ�{\`�?�|�4�k_��~���	�����gQ569a�k�R�/$_e�~������z�PN|]�&ȋ*:n/�.�t-���	�V�H%�|�F��.�w�I��_�N4j�v��A~?���r/#�ل<�Ss�a:�)�U�,��ҵs~u���n�__h�|ðקQ��&f�¾��'0����G��7��X	��t��v�B�������k�<D/
/�Ovn>u~\zT���[�Z�h��	
���Mj�",h�����r��sUT5\�mU�f>[� �H`	؂�_���?��0�S�s|�J���ܹT���S��f!�[vKSR$.i'�J�\>=k%��Ծ;�N��I�1+�*�{3��q��evM~�a��W���& Dӳ�RB�<-�ܨ����0rۄrqPW�yxWL�r�)h��������h3����\nqUs	��#LE��!��&+�ޜܙ�3���|B��N�-''jd�q�D�YI%Q���������=�y�������B�����L����
�� ��K����'$��oe��w%�'� `Y8�zG�z~��qX^汥���[8~ƫ���_�}���,�װ�.�U�@Aŕ�d�Ԗ�6�������K��dN?��ͽBy[,������"=��Rx<��_�����8�m^_h��8���)�[7/4�R�N"'!.�x��n�3a}����5���D�M�(TP�X�Sf\8�B�A��hq��;�@ώ��������m�8ouy9o,aɇ���'�)dkɼ��R���m9�Q �}�oFˀQ����<Sά̻n<��'讉����0�0�H�����`�>�>�� ǘ�p�Y��oX��'�ȂCG�(��l>����f̃�XFno2�q�ޑ���t[�9�?�0@�"�
I���%���M�(K�Ƚ��qtߣO(�Nh�������)�Z����^s,U�Q��6i[�M`"Ϛ,��Z�ؑG[�[���&v���k�����8�%rRވ҅���iZyd���l�z��|�
�{9�����w���R�S��YL���:q�6)0�ù=�V��������=��rH@�(	!��}�������mߠ��2u���*�%�&��x>�~Q��o,r�Y���E�'��ئpb��"pM8Y$�uҊA���2�i~yBg6!�Nk�{=j}y������N�T/a��ċ�91������:�B2�1*A��x� �zF"Mi���R��I?Oഠ��ܖ-h���fRK�����ʓ���݄��~(�C��]����kk��*��]Q	r���"j\J�9ݼF)���x��V���攚�)��-���湈]{\�Z�����7Hk�Ԓ��aܡ�z����d��� �W*�NZ�yr�0�_5ߑ6�;� 5��;��'�π��i��Z�H�ɰmK�C����rE��R����>����L�$�&���p��rI^�4H+e�K٥���������� S�����
�����Y��`%�,�
���Q��I�'����:��HP& ƢrR��0�1K�b�Y�ݯ��'�DPJZ�f6�c����q母�u@q������r��*�0���6�x�y��.���ވ|~�Z5��h��
̒�\׫.�l+�[HͶ$5J�oF2'bT1�&|l(.�irxkz��zD�_�,��S;̅�aƄ����k.n���Q�6R��y0�0�ȩ�>��J�yG�H���%4n-�sk]�3�Jyg����י��z�h�vE1B��	^��efп��\\�����"4���\�̈́���9���/�i��m�M%���E��i���ϒ�����/H"ҟb��T�%48^[70oEx&u_Ď�Y��x5�-91kSY�@M�T_x�j��]��S�xvy�͑)��gZ:U�A �Aw*�����R�VK��1R@�p6�lo8��8b�UOEn���1cTl/�d �G�����R�j4���N��o|R����6�Cx�,F�&�nk�<%�ka�y+��i� \����*~�a�8m
��3RJ��G{���������v��?������,ȷf/�k���υг�e��L$�������k��Ӣ��*�ɳ�B�@~���Èru�i���Z&���BsUU��P=
���|]��U3�Q����W:r�?/�!b��i��A^.�1'=���?)�DM9����K�2KQ�p<˶0'��/}-S=�eƏ�!E�(���W����+�5�e�S�͑?�^#T��0�H�w>Q��'�}ޜ&�F7������Fw���y���5�&�G(��,^�dM$��_1������1=��Z]���4B��g�iS���Y��1L���z�um�E�q�ժ��ڻ��ZCEÎOq�' �/m��<$�N�.g�dǤ�@\(��a2QS��\�]s�GEaK%�I��^?��^
���L��0_O)�����W�Mj�צG<�lzD�x��7����Z�\J�J��=Y��Õ=���	�M�J�7���o� ��8/�>�j��#�F'rƇ����,,�P��H�i@ޥy9��S��/J����<��5M[P���U�P��䛱^9�56J/#V��"�(�ױ� �^��4��3���� c6��Ukǲr ��!񙼹d�Ϲ�n�4�,���� lse\19�����9K��|�2�!r�ֹ$?$�4��AK�-ۚ|4���B��Ɉ���ȝYŹ�����T!�<��l]��F��R\p�}}�$���n.n0���B8����6���)�:6����LmpC��c�}}��mF�dS�������o��=�U老g~s��r�3��FE�
�΢}usc�{m��h��Q��i�q��q]��L��nn�~��lMrW]��B�ozUZ>o�$��E}�%��>O0q&~J��.��ѧ� �´�!��1g�@�0,[r�4��\L�#��$���F�c�l���P3�\����|T�텐_����̞�G��E��S��X�:j�LW���慮l�'V��\�S�V�̣,�����Ձ��k
�"��m�rt�U���a��W@�����[]�уS35��Ii~��!m4���A��	[���d��	�_�l����w=�Hh�U�s���Vn��Cr�"ΊLoУ^"l�|�����+�P�"9d��� a���k�Y��fx�yy��q�y���{�ҏB��91�	Z[^�P�*5�DS��>z5�}�9*ӈwٷM$S��l�i�}&��>mwX<G�Z�S@!��泝�Qg�9�/��?�]������$����ʲ͞��`{��������n��a�{x<~W��9��M�hĿh�9׷~���	)>S�P�Y��\��WL}t;ŋ�
F��a���$&Ⱒ�򛌯8���yMn�2��YNC'�殐�3��伔(p ��؇��>AC0�X�ȃ�!���̌�U��r�a/j&����|jq,V���n���Q�������G#�"��2�vA��	�Ȩ��v�2�j�b�?�0�����D�M8�4u�����{J`�.�_n~Ba�oA@X+ջ~����>^#v)�7Q pD�	���A���wk �,�[:T�}���o�A(
�7z�$��D֦�]���{�I�$v�괅�a�����U�X�me���bWi�pB��%@���\���n��V`ѧ�����Ɩ�?Z.p Go��5�pN��ץ��1�d(����3)�m�"I�cp
���2�L#�1j�"��o��[�^G��Ч��0[�X�^�
�.`����d`�Va�V�Rf�*��ªS�`�Ҽ3�F�zhy��m�J��$*�y�G����h�u���{	3�T(77��ų�TNג:G�own���^KF��	�%��	�M5&��r�?H�9^G��:w��"/Z`f���5�v�ӹܺ�t��(�@G7x� n���e�5�\�Z>� N�8��6�����s)�%*suһ�|��(aw���L�X�3A���u�����O�m���o:f"�5^���M�Է4��Jy�l����H�J>�[�k�үT�H�~ŵ��(��H?�h��/�f�Ջ�n�\�I��+�=�����R��"w�{�i4��J�KO�ѹ�õxs(,('d*6_I�@l�n8�6�6\�M�'�W����	^�	�f��/klb/�%A���<�{�����˖�d����N���(��r��C�6�Nv�������Qt*uf���ƁX(uwA��[�ϼ=$JR�3��9��3�2Vf��v�8N1����氽�A�5��u�O�4a� D1T~���O�&)H%g��@ైwJ�E-�R�D������������4��$���z�빙��b%C�n�a-�fן�G�]�G"�+X�k��H����Uq��B�v;P)��ġ�Q姼�^��p!��rm=^ؿx6���Ó�V1 F-�0l�iv�A�ɦH�IN��7y�PSi7�ê��!2z�(UA>��Q%��C���g8��L�.�'��"��^gFe������"#|S!��C0��;H]�X��4)����+�2w�y\��$�2E��|�#���D�M{�.�5�P��Q��l�~QJ�}.�'g_���B=	P g�K�K��������2�H�|���(�Ql术cr�<��#D�t��CiI��_�S���
C�a��ߐ�n%K��4��~�f���6we�,���09>߀�:,ƣG$�ZE����P�=��|���V-m��`��Ǖ$�k0����(�Ǖ	�	�0쏾�͕H ������˻l:�m b�B�����K��l@'�������1����!�+�������5-�]��d�%�zz9���א	�+óīX��=�	��R��ѭ.�Lp`�̢3�H7��q�&�Q`؇�V�y̙��|�s��)D:Y� �	��r�
s@OeWp��W��p����=�H�2G/��E�B���M}`�ˣpϔz�*D�t6�4�[�^E�<��� WWs1�8F��梑x ŷ��W3�M��іg�KFh��sG`�W�!Z-�Ǔ��n�ʲSj1���{Ī���p��t��H���	S�+��'�j_WG{���a����������K��f[ޝ2�-�m$�P̧
��y�u(b/
?:@���T+m5��w�3���u�7��W;�ĕ[�R�#��JL0��)r��3�$3`l���^�.hM�6������ʲ)����(���h�Uir�D�������!+� ���'�K��^��D�C�	j#�7+�b�H�<���չ��6�3;�1���z�(�����{v�>#�J��'O��F+�(�S��͂:b{ܯ��L��	}��ޮ�Ĉ��b�\��<���|���
sg�߶ـ*�e�Wu����#ۆ:r2<!F�Q=2��AΓ��)tZ�~�V�b[���-��A�Z�<)V�lr)F�� 4c���C�4o9��*��T�\�u�\*�'տس�2��v"/�~�'��>$�b�m[�`׮��A�0��OZa����Ze���A�(AS��������asV;�,%s�uU�J��f ��]h\�B�׾ ib��4�.�Ƣ�	����Bkˣ��X�Ǣ&�Ul������'qC�c�TV�>�</@����G5&�e��1g�"�m��_�+�R��?�_������Ϝ_P�[�(e��(�����tRڢ[:ٕ�GEAUc��rс rO������5�j��E=�7�y.m�A�C��]���H�i���V��W��]c�Rj��&1>:&zc�PWLG ��S5�}����F4��GV+���,EI,���r�c�!��z��4��Ÿ�/�-�yA�E���XaՈ�ޯ��E-G_�J$}
��|A��3^ևf�O&�yL��S�ڤ@�	����4:*50M'��<��MCD�2)�w�����pK��v4PFL��(��y��o[t9�v��Qw|�َ��0����'!�.�w+�%�ֻ%����_kCS�����\)���-����HQ�����r�SL�x�:�u3K� y�c;~ѓ(?����#֑���ʿC�:1m>�k����Y������$ZA66>'h�k�w��U8%" Y��h� �"���?ܘ��s�5S����X�aAr������o�� Ept|��է#ͦC��zґ���7Rʳ��h�p���(����/x2R��3��	:�v���1V�p^j�u�F��We�W��Md{��3Y�!r�V����'5��_����B��"��R�\ ��>�T7FNr1a���2S�j�R���̘s'gL�Q�>��9p����6��e����?��Ach	��0x�d�v�.�T�8���RT��5���T(lF��wK���}�����}HF�&K�vj��
���~���١��PM��:{��6!�Tc���84f� �4���^c܍ߙ1Atdv�:�1����,64��Ɯ0Unm��!.S<�^�&��tZ�-E�eߤ<ش[lم��Ln8��ӆXE�Mv��+�dÇ������Bu:�tq��ǥlw1.��3jH*�+�+��_д��}���Q��1�B*u���F!�O��+a�J��Ǽ[c~x���>�A���4�;�>Ȥ�a�H��.k����r��!8�i&X�8�*�0�������Z)��A��^�j�U��4���j$�6�u2BBL�C�S5R҆8��*�r�Z��mΔ��b��ݹ tY"����9I�h(�.CH��c���ƈ����w����5������`J��F+B�����ٳ�����@mr����uB&��l�U���Zk�I��.��l�0_�<��q[C��`Jd�:����"��v��+�t�p�`��l��pE��8�C��Ռ�����^� rnƔt���c�uh�vXp+lǻ2�֑bc�2��c�搢 �m�ԖOb㺴铝�����Ij������L�����.>�TyЛ�(���h�)?��.Q���lAi��	����J7�e�J�X����$�u��o�z��G?���ZK��]ʗ�K~���ʻ�kEB�AF�ۆ+�{[k�
���re9�LWA��F�[����w�W���u&.��B�dV�4��D��v�9Go�)�zx��U	_)ؿT��E��v�̤쐗��AF�A�"a�)T��F�7�5K�P�e�����L�{��K�vaW�N�16(G@&:��t���@�M�e&�Z��\�<�������A�G��p[��;Q� ,٥��"e��Վ%��rw"a��s}p�3y�e*��5�,ı��Zx��ud
l�)@�P}w(�`�D����3��6�+��0u ��@X��M�_�zx Ey�$�j<4'P����k�d�X?�фAD�}�n�л*�����0�#7���b_�P3J k��Y{Q�����b�@~��٨�]/�?/Y��g�Xgڔ+@9�'���(ʒ�^�݉��C�a��ʭ8���w���)��j�*l�ئt�����S�OT�N�;=���G����]�g�v�7��QZ��-ܠ��r����.OmY��¿,[GM���t�$�] ��/Z��[��Ҩ��8�u)U����/K�:`��&�o�W���8�X|⃉���ʰv�o�>0�y�K���b;���uȟ9\�Wc(g>��ST?`d�w^h�{{�q�{.�;�9Ĩ݂�~X�bHN�\9���:%���4�����[>,N�n~K�ZQ��^84cl�Ш�_�Z�:�w5~�?�Ķ�f �{e����f�z�`%����<�:1u�q}���b	����ʧ���#���\���!�&�}�� �ƛu��&�j+�Y��+�}�f���D�V���@F�`��=�ؼ�������~��,g�~N�����Y��B7$W����S����:���	}�3�eJAl��܎��J�bl#ЪO�:���k�?������N��A%Ș������'�	}��q_�������z���6��g�WU0��k偦�i�����AP��!r\�9�� ��ع|�t�V=�g��|��R9�':�K`r�A��N�F=�S�U(�b��p��b�qi�D���'�*�td��4fcߟ��"_ S"���\w�!p�/�_Ĥ�y�T����)1��3 kC��n�kז��4�Ct鷕BCE�� /U��K����HW�2a{�]�h06�{�m�� ��qH�I��;T*@��"��E� g�b��[ r� KI-9����;�y:�&G�e��!��Q͔�-t Ƀ��)�3��R�G�"d�mq5p��M�.V�@�;�'�)> l%�E�CӦ���|�7>����x�������� s�}����ߊ�1�V��#B��Ed�<%+�UJhS�Yfwb/7'��҇0d��"^B��ݩD�ŭ	�6N�HH�u�T�(\X��� ���#�2J�T缺�
�'�Oj,;�&�{��&�z:@�#I�x��OQBO���N���Ϡ�i�����!����r%��k�_���С���s��|h����=�������wk�F���������b�?}nk� �z=�d�@��������1�,�?d3�NNZ��w�W�I�n�<���DQ������V���	���}�Z�l��}͞�&EM�]�FH�'�`1p��٤ �rKk4}���5GM`�P��?�0�޻��^�b]�#F���?�"n[�䏹�c�s$��P��x��P�� T-��[4浑�P���@���v0�i�U(s�U�X���^}�Q�zy��x#U��k4y��-�	�U���2�O~�`�?�+y���:Ŭ��4.�'���尵���;;���s6��="<7�Lv,;e�ՆxJ� &C���V�e�
��*�f�	����y�2�k�c$��2�Mt���=n��������Q*s�M��#��t��2%���o����i,��
��h�ض9�Fpo�6�eX�f���N�[�L��^
R�O���G���)���Y�+�쐻��y;���3�*�|����-��Ic�BO�����p�Gz���4R#1�-�9SZ��W]o�LG,�h�I.;���N�<P�kݾ�R�R2~��w�����5�2�q�]�)�N �1�9�⾋o����o���z�N퍂�bʹ�gE���}^l�ٛ��\J	:p�?�g���nn`�hp�Ȅ�#�	�~I��-h_1.kJ�f��

����;o�����L�1ء~�l����Tv �4��}��[���zhL74��� ����>�,�f�K󺫨e0݇�C���gӌs �i�=r�Z�$[��=���0����ֿM�w��̴��>�E�u$+�[�~�6հ� �'lzWy��`�p6bvۉ��O*��e�9���R5�c����Is��װ!�|����A�,�G��&2�l0۴ ��T�ͦGD�������P��mP����ᡌ���]�������U��;�L�)�i���d�"��g!׀����\zG��z@�P��������_�f�ϧ�9|��N��%o�8�]R�w�^��*��ڔc�!iS�ߤL�D#�gH�g-���y��!�����V7�*b���dl������20(i/|��;_O���T*~T�)�{8��ԧֲs�)��J��,���.�?{�T5�^�3r.BZ���C�˘ ��=(��
ί=�TE#�/Q.5���~�ۜٚ+��4�qGψ�y��1]�+�����7�mA/'�/g���Q�l)�M���c��b�śo�������h/u�Q�4��2�id�f�[�K��5��Q�[�٩��`_��E9ݛ�'�]����>��[�x�c RQ�;X�����np����`2�� �zЫ�֫B哔�sA��Ld�ܷ��G�04��$b"�]{�K�D��o2��
�����f!T<z�Gժ&L�)��.]Η��ff݄��΋&�BM�:V�*dB��xe�Y&��`��� �O�i�/uFN�~��L��l�N�.�]d�i��4��?kY�	���KY՚�v��Kc�)�G���-�� �GO������f& �(�L͋
��?E����k��5>>�i��YAG��p*�;�kd8�����=ufp]*~6���P%�f�խ�Z0���^��)�[Kj�8\�hv}Ĕ����?�[t_ڒE:�Ɣ��F�a���F�~����J|v�<u�P�����Bv�lG-�=ƒ2�0��&c1��1����-1t�S\�r�^걊�t�]���o����کق�w u�Px�kE�����|x(G'o,��T��:p��<_��8���b#�_���#���C��h�7q��j:/���\?�y�H�z�u_C@^�i�z	\�����?5��Oa6q>ҏ�ݿ1N�I����2k^�-�NXOЂL�����h�h�GC�񛩍�v]o��B�x��`�mx^���'��G����0֪�����A(����7�M����1�p2
����ӕ�.�L��j���/qKڿ�4�����c�x���^ǞÍ�j�=z1O^.�^iLG��]��
��p�Y�]�5� {kU�5�8+�0�ʊb0Ӌ(�n@��\�-�#�^|���y2֣�I���`��ii�褖x-l��R�����y�$�t"�4{l�h�"���v�3���5a�8�Ef���e=��sg�Bm�p$ �#���Blz��J5ѭ�*͍�e��R-"h�����}�%w�')%���y��X����Ī��eI�I}F@#XE����;	�Ui�����o���w�w� |ɠ��f�C�q*j�� ���1t�a<	��~^x������I�6��2 �[��$�À
�o�Q�9��|�+5?�e�u�6+Gg������!��İ"��z��n�F&���k�!�&t�OvmE׾�_d���	_���i5�g9��\�g<�ORk4��@����勁���g�-t����{!'�c8�z�X���Y'L �MU�����5*��z���~�#�,��%=2u�m�v
2	y�.=|��#���{�jȥRN=�X;����U�b���K�Wg7��5*���Eb�D:����R��K�������#��P~o������u��0����x���3
$oBE���ٷ
���	]�7�bHj�hQr�z���R��{�l2��� �,^�-�זK���}s3�J�;l���B5Ǫ3~c��؟�nDQ��n�0���/e�d�d�"�	Q�R��n�ր"�0FطP�d�.�r&X�3���x7��;o�ц��,��X��g1�q"��U�(,���Μ�Ap]p,|4{� �L�2v0��]t� ba�3�8�u�`�ZԚ���,Ж���:��ǽ��<a(Ւf1�^N����H{��oЍ��ys�E���6׸j�����N,i�v��+6?��^���\�)0��x4�-�DN+"*��ճ�E,3�P�z��w�$�}q�d/80
n���U���zn�D�Tv��n��U��v�kb�%F�0K��<m�$�7[�����q`�=��k��ʂ5��h�y_m��%��g��>!�AjD3F�I����27	:N�txQS�i��}�hL&Z��u� �Y�7QӘ�7Xv��}�J<FE�l�FK P�{M��8��b�!���%���3J:��O %06	!E�ч���	wkI��P�.z���3�l���������'�hマ9\q��+ ֿ��r�N��m��k��X)ׅ:*��?����ABqXJ�Em�NN��q`�+�	�K�-�!*^��PzU�&��#ć�i/��O�J\t�L���(�������E[��Kq8
iYs��A�B���Sf����F��R�����˅�@��As�^[��V����`W��W�|��B|�.�_�̩5���������0kp0p�"�wE�+/����7vo��o<	��(��L�O��^��Αqui�f�w�XUXR�aM�2c�X���4������:{Ȅ�S9�V�mU���s���X�J��
5��À��4/GN���v��[ Mi�HˢW�oB�}8�N8~�c�`R�$�Ku��L.�
~YYUۡ�ޣ�j~�?e�޴P^HV!�~ذo�b�O oV����47���Mn���J�k��X��?��Y������e_��!�ݓ��@�&N��N8�����%'�9�W|E�$�|E�Qf�v19�jvz��i�l��,8vQ�3|6�7��߾g�o5;�I|W��x���H��<�+�G��*����t0:�ʍq�>k�{.Hn͹� ��R
w8"^ ��;U���L�ɠf��me��{�)�����R�����5Dt�Ӊ"�%���hW_TU�]�6wyt*	�c����Ѓ�x�`cZڪyT�+nd� }���8Ƒib�˽�l�̥�Ԝ��ٶ�o�)��U_�~#�7�.#N3��vx�l"l�)b��$r�v�xcb�6�����% v�5iy3!�5z����<A����+���k5��50;I�*;�5�@x�����1W����m"���}�+��*���K�=I2��)oI����mP�a*`��x����z��ӀV5)g$+���/Zc'�dM�E�%ݶl;��!鴚�V�y�u�+A�L��j��h}uY�+��3���	��Y�Ӱ��=��H.nKvUl�@���?�HR��E�x �d�g	�
Cn�9���G$U����|�`�y��t!��٦B�p���јY��z�ѼνK�
� ��d��=&��Km$EL�׵8���D��I�y�^��6�����3<�`�r�������zm�!3�sU�{���Z%`�R������x�c��@�2��-o'���%�ϥ$�rz,����i��@77)�h�vP�O᩟z��H]n���0
 �ؑc��Q7�"]."{؄򉝚�7�ΗéS\W��J-8� ��֥�%������>
_~Q#���9=�)�ј��Z!D�W�\��5�=���i��E*�~���P�:�v�T
c@?t?3!q�#�}N�	���?p��1��4l$�����bq�1#w�,J\6OS�������i�ʈ���_�Y�b�ꆴe{��U#�S�2I��~A��է��6�V�(�&���_{��4 �������R>�o���+�cҞ~�@HIq�7Z�ʶ�/V���]J�U@��~wx�K�Xd7{^_Œ����6��,��N���U�����@1
P[W�M����3�Ti��?r�(��.�@8�]��8%�c޷Z��$ӹ�/���
�_G�du�(�*�HU�M٭F�ك���*d�#m�ۨ����i<`��C#A��2��
��ճ"&n|-E,����7^=`.�~�;�Ζ�8�e�Kԓ2p9D�����T��y�����M�����B!�c10�0A�*�&b��87�g�M��39�

���0��7�+��q� ��6�fG������0Ĵ[?,���i���r��q�h�0Δ�:�dV+<�H}������1�qoWg ӵФ��u����Ɨ�·yz�s?�n}���.���;�j�5�������FNJ!�R��r�G<w�/K��lx]�7���E�%*P�ޣ#�D=�L�SI6u�U�0�wH�{�����n ��$�_�q�p=9�1���Fԏ~"�%�ҹd����F����}ρ.�r�`�Y������l��twҶ;�s�s_ld�\O�O�v��k�t�x�6N��e{`D6�'��[��5$�]kQ㙚|��;v��A`�⯫mu��>�c��:�D�!JtH�����]8Lr���}B�"_��9�{@Ͻ�E5\��z���ve_,BF?A_��&�U^�8i`��
w���-�^�9%X�q�]e�dJ��zd'O7�|���IO��9���V'��zN��phB,~��#�d��o�Q(���i����ڒ�f����V��&he���_c +q6��R��ʹ�c�7���'v&�!Y94zQ�0X�~ޠ���gg��({��JWJ��o��3w�0�e�~��L۔ N��קi�Y[����/��,A��q�~h��-d�{͵l�O�1���X�e�����m����Z���C�<` �^G���\����Q��w�CϖEUN�Z�u�=��ѭP<�(Ӏ�h��S�
R٨u�(��(0T�P�#�ک@�̮MWK	�%��i#��<�Z?���bӧ�yo��-�[�9M���%��ͯ[�=�� ��q�*�����~�1C[ bx��,���(�+�*�ٮڗ�JJ� ����T��丕8
wKw>?]��Z��{�6G�j�ȡ%v�*�qe�-��5Q��O�Y����L�*��5q������i�d}���9���;�s������ĦdH]��S3��:�f`�);�x���4���a�]o����z����$���^��� �
y�J�
G��xr�8��ØBbEA+�r��g���>�b0�dlb��[bp��j{�_�{nE}|�'�9�nG��3a�b�~���3q-ȥnx�����;�_k&ƽ	����s'�u��]k�k�u(��5�ܱWy1��
��
I��x�m,��ࠄM�]k�����(�As㬶>���_��z��9V�>�Vzc��A�s#���	H�xl��6-�7ń]�G���~c�� Og-��y�f?�g��-i�.-��|>��* P	5�*G�.%"�����8�͈���8�k�c eآKQY:hB+2���N���ծOX"�{��C6�g�3��a�� Ak>c���ha:��>K=�3�����b	3���B��A�HA��3Fny� ;�N���<��'z���V�$�����R?�I�D$�����9�ɩ���ݱej]�d׽cV �}��
ȚQ�C^��V֢!�P?au��jD�f�Uk��熂Uf��q�5/b<�ʏ=��'��|MH	LTmx2qZ	#2^=��6���<��~�m�~לּl�`~��`r����C���{j�uzv�q�����+7Q��u'K��xVx�`7 �E)��Z��@�S�8�bC��J�ra0�Y۶���ۤ��OY�!T�-u����Z��P��Gc�K���|�߳��|�A7�Y?*ߗ�?��S��8I�){W��aX�5���]�(DW5���}�y����r�*�r����֝0e(�Y�7ۓ����������G�ș9�\_-�w��0�܉r	Rd�({��-
,�{�ؙ�Ť	��؅���mJ0E����b��>o��������t=h5��T�]���v�O��U����N{kM�H�p�o��2�)0s2QF�*q��0%����.c)�\-M���B��᳃��U ��c�t�H�B#�d�;�G4���tO���ix�
٥�5�-�S�/e�V�D;d�c��e�V&a��[&�������� �=W��?1��o&�g�t��#ё��VB��_��vFw6r��Ev�i%��C_�x�~��ȫ�/X�F�RW�6����`b���']���/����{�J�ݝ�3�ʏ"���y��#ȍ��ϴ�F)��!�.u��
�g��qf�+ђ�؁����N3'E.ZC��>w�=׊���6�ԩ�����8���sr�5ժ�T�fюK��&��b]�ͣT��b���8�2�!3N�7#���GwйZrS�8�h��L��#�`��?�z�r��'B?�ow!a���?�ǃ T�Y�U�%-3-�.�K��j�[�����0��B$�]�Ф�UT�g���;OUt)�5�l.;kI�O���r��M`�Sq��foh5�o��d�1E�5��j�B��Tp^S��e0����0�u����a�Z3����:��J�E�04w���-�{���cd�i?|�|�G]� �}��^|�dg�B�/����n�Q߽c���=E�W����{���M������/�z��%�L0�L�2��KǹJ���tX7g6��Hz�Ӊ���؞�OJT�f��;y���5���E����~) *����������t}�&��B*�.�R�H����m[˿oh�U�gM���cl�-Rz[�cL��M���;�D��RSY�ij>�8��E��L���L�\�R;3�W�S{�,�&z*���n0N`�dщ�fg�wFz�fއ1�c�q�hTa-��gK��_�̛�iO�3��a3������lK��:�c؛A.�m�l����8�pST]� +(~�҃~��r��*�,ׁ��W���v5�8������e�8�;B�����yx�y��ٞ�N+�PT�%��w�c*� ��v@�ۑ~AFw�� �+�2���dk��bA���F'C�h H"���Ru��D'��P�/��,����$ì�6�8�e矚�^9�X��ə+j�P����yJ���j�~T����֨�~Л�v|�F�V�a���7�T� G���S�`Q�@�V1��i"�3�	5�M�a�)$T�����&���T<�@N
`��#��Rɷ��c���"#���.*۱`|�N�@�k�r7�k�^O��D�j%RuĲJ�/��s���bw�L����qnKPM�UX���q��Y����0*9��. J}��� �̫y
D�T}���i��kq�Q���ٽ��j��r �)���Q��WC}�C�ְ��o��.Ka�t��x�w`��x�]��'H�cTM�&W$��q-�$��҅�?XbŹ7���7x랇C_�����l����9
$(�)v���fV*QƂ�+mG�H��C)��G�b	>$��b�ߪcцk{��0�A�)d$Z�ۅ�n:9�	���m���K�cL�۷38�E�&ϛb�	����)m�g&��q����J�u��î�f!��
������p.��:)/�P­�E���qdW�B��c�c�::�Y����H4������q�.�75��E��+�>��?�,xu2XY`�Z�q
�����
�1�qb����頍]��z_��p:��o���Za���5�Lx`A?��ꌚn:�(�"�s��.�����a�-Q;2�#t�2��\ĒH���d���B�K(��K�b�b��3x��V�m�bL&ՖR����Ud�̪A3�!����S�P��d�"xn��X�v��Nշ��ߺ���]f`|�<�i��J��֡��-��\W'T�i&St*w�ZC�;�) �C� f��@�n�E��ʚN���U lY�9���΅���^χɶ�*�;6>��R8�j�{���^Q�8�F4�K������^�O�_���٘P��G#��:Bo���� �J�f���.{���`YX�0|iL�<��o��h�n�^����q]�Q����� L��?�G�KiQ�x����5=�]Z��o=ě��?x2����A��q���Q��!4DV��ѹp���@5�m���+!or���?���b>�tg� ��>M��$@Ⅰ��2��
�U��b@ԟH��pu |5�"\�pؓ��@��8	��_�,��h����� L����IF���$t�8��U��$�� ����R��[L=�����*ʹ{rؕR. 5��7�E�'�Q����	igg�@����D�
��-7��ڕLn����ki��u_+0_�P�����PVZ�xϭd�m�'�^��J!�-�w���VB��f��x�:�&���P�����M�1f�+�K����5��Ai;H�T�Yp�Q�䔁(�x�>B���JO�?�t��1S	j�%�`�A�����na>?�w���Ę��;�X7=_+����.߂Å�;�3%_�k��y,�i�'Λ�b�2�d��3_�[���~k����=�x�ȁa��c�b\	�٦EEҵ�@ O\����O�tƊ���E��{��7�l���ܳ;�.��^�y�rm�:}�f�i�7�u��5AJ�f�?��hUy��17�J_[��.�/��vL(����Q=n���:x��-�	��NN���n�>|c��Lڜ=�����Ac�%���Em�w`�EŞ;1:��܄4���(����w�'�QER���zk��|Ts�SfW��f]0N�O�>V��d�(�iߨ��N��噉�2"l�
by��!�R��^
�b�r�-$?�CtF�_!�y$���bjv(8�� ��1�T��i�Da6\��o:l��v��vD�[{����~\�>i�,�|��a�5�(#�ɚ�z1��h*9N��^�ۭ�;^��`u9]���$��4&O�׍"����01��H����gK��L�7��4������񪮎���X���_��|Ch�~K�"?8�<g���>�m�-�"V���9d��D@��� oI�7����r���9C���I�@]�2���"�d
���Y²�Ҏ~��0�g��cp[\�WZ!�}y�+�8�\R�A���z'���9X��Q5R���t�x�1��`Ī��m�����lkԍ��rB���${��!���"��<����,A�������bѭ��(��2�<��l��������cNA!���ڸ��op�܅�эj0�����U��\2�2�~�F5^*�.��۞a��y��L��)��L�V�;'Y���C��4����J*<��M1�e�{D�-����OPW��[#'�pu�	�o�.ұ�)\/���dF����G�f��`��f�j��|k�E���#S��q�n�6'�e,H��R��W��j�h&0q����햼k�ܙ�_�
���!n0k3)E��X���(6�]qa�?����%�w! ��{�C��J���(�i��
+?u8��(+ZX�-��Ȳ%�����>�p���+ю)��\���{dA+����s]�����CV}P�Ľ��[�-Ry��1g7�qRLI3{���J�J���$#2�SY�l��֗��#�vx��Z�Y�{*�����`��F*cF�*�6���D�77���JH�zV��/�u ��@����%�LKK	��V�84���ϖ;��O`B�'/��EGa��a�x]�rm�[�[J8�}EA�kM���f�9�8 rx����Sv�_5�$�tӘ����Fd$=�-�Z��@�_�7�~߭�r�	�ݥ ���OD	��`hJ��L�f�I�����8��f�꒮� �,Ζ��wCL�3��_DV�v��2<�Q!A@!��cR*>�h i�>f�a�8�"cq�cagޕUd5m�߶��g?��_��*�]ݖ�����ܣ���='T�q��ơ+�� ��ЏI�Qh�� �E�6�K�aw��U��u��O�?�� g�噋�5��@DPM�6�|�t=�`�ɃX�ɹ&��}�/g���-��@�D1�>�,vY�����
ה�:Pp=�"�cJ<��a�ӽ��ʎS@t�3r�ˡ�3���A㷱җQ�{���W�`�A���߭~0եⷾ��z��󈍶����3d��,��xe팂��s���T�V��I�s�g�����~�_sE�����1-�P��-�ۡ�\h|�YMg�-n�A͆�a�V�a���!xB��t�� Js3�㕄.��I�Jh+�cg�x��.�P�7H�a�^�!B�(�]��v�[�ь�4����wQ
/NT�`��t?h�ݦ�^�ͣ�ˌ � #����1�X��D� ��,�Q8����T��A\�GQ�?)�����5Haթn���������	/�[5�7b^S'KDs
�����^MVţ�U"�\�c(����;��|�|.�9�8ؒ@] jA�+�r��(4�5�t�L��`�1;qXc"�f�������W��&��|�*�T"0�R����p�����]�f]K��N��6ǫ:���>SP�P�'D���M6�:5��I[���q��=�?�����А��\�4Ռ�S��=d]�a��P!c�;��I!�B�tB&G����D��8ziS�`�����l�"�=Y��sl%�����+ z����'E�bȬ��`F�|�~��s'��B�<�#��}�̺�Y��hx�5�j��}��_h�C}�Xi��2����i���4�1�\i+�i=�������D���&�;~w"T�e��%O&C�n$!�Y�i���\_���+�[v� ���p��VU��(���z����ڷ��!��3ON��i�=SDBt��R��+�y��wM�=��J�|���	��aź�M��%�^N��E�ŝp�L+,��:hAn�[�)����H�H�21�/�A&kY��B���Gq��#��,��7(��ߞц/ �M�	\�r�ӢS��}8��2d��� �+�l�,be�\ê����.�T�����hf�[� v��I��?x�kd����4$��<���Yeh
��i���1���ͬ���A���&��Y��;"����ۻ,�$��������c��2#��H��l<�����{�2*�z��);{��4e&�\���5��^��@WYzS�Y���1�e�ډ��2`�Z^�?��m�.�x�>��3M�m�|M$Í�k������i���p��n?j�3�d�~Z~q:�ĒzB7�4n$�He�ăAP4�TDQ����on�M=j1���t^ls�{�V]��g���뾭�7"p|!���j���i��|�de[����db�c�O��a������b��[~��E�w龎ŉ\�������o�'ɈcE���?}�����/&I��w��\h_�u��n!�Pa�_�y^c��X�Tk����yg��.i���ΊioV�\�v)�G\śJ.	��<=�_��F���>����Y�֛�aݐ��U��f�/�c��xc�ſ�ݞ�h�l)*%y \š��r��s��m䙋�$)AYBl�x!�
χ=e�:��"(r\�Y����!��>� #
�9Қ��P���kC$�(��&W����(r�B�~�>����K���U����&�[��_����� n�#�Ӌ������̶.�*��>��$����|,PC��6)���X|,2`k���|oI��ӟ$j���w���JmRr?�Z�H*����U���ʥ� F,�k�Qp���:�:�:`�@w�宾��~��$�Ծ�F�*�`3�����Z�3byL{<�G�r��2
���;�!E��p��W��V����H��+ӊ8\��͛��Smf�)��$S��+N`_�M[)�>B�|kO:D^�Fʺ�Oq^z�E�n#խ�Y(�9��q���E8<%ʉ�o�l��L�G��<����q�06bFI��K�1�IP�ʞmާmm$����3Q�Y.J͗�p�AyS0`������ #f��t�L��¨t�"�E�恊��:7 f7�F�I�O����ʚ��ݥ�,Z��?f���%�-��iU�=�+�m�ݿR��4�'�jˊ�T{�ik�7�9:��8�ɺ��*}�T�F�>�<b潟&�uO��7{e��I��=�����4�N*�y�@���46מ����[�׵��-u�s�
'�}�r �[�?c�L'�Q*1�.ڿИ���>�������cH���F=���>���=&�5IJ������>�!`�2k�:�n�vh3���/߄ԥ���P�	�n��N2�(_hkݺ�u{~�`<gS(�`����e�[�1\��+5��ES[��T6F?�~�0+1[r�̍���y/����w�r�±�<1����o
�颂�Ǐ�@�D����
��W+-��9�TtXFoS+�C��ף�f�l)�P�u�q�(��z�aPSd�2�~���g��DC���d��������wa(Ę�����K-���#�"P(���*\��`��*:����S^��\O_���*����Z֨��5 �Q�1����ƶ��PG�:ŉ�;/�$�f�˺k�/�tM�]����k�!U��Q\�t�b��3�u�y�{8B��Tܡv/#�ҰO%� �A_�D�P�}`��kS�����8K��/0�'�'��H�;*�rs/�&�LA���2�k?�w���s��]�hC~�`;��2qd}���o������t�U�AԮ	^6_�Ket�~��^"K��_̞$�\_���ɝ_7ʕ�&� =������p{� 	��(76"7��ۏ�%�0��@8�g�����V�ϋ���gOw�yQ�����Q�%�UWy�;��l�ڻ�Q��	@�F�O䀉��\�	����цn��UV=���d�H�	���Ƃ�t��2���!����:����Jc�<R��4K�`��J�N���
���%�TV�� C�E577ы������s�p9�
`����a+OB�(�?������ߗ��MS�b*���VK�:�\�o��%9�nF�4�gl0��c�p�9��O-�+
2��kG�0<�#&����;��}��:q�S�\o]�Ȫߴ�T=�%f���ԃ�;?v9zv��Lf�
��9��*J]��$M3.���j��_7������ג�������k��Q����d͵'�O��.~�U�~��M���^��'	yёQ�D"���)J*�74�|M���Oc�]��*=���ᙅ��ݖ�Ը��� '�w�!�E[��d�]�#�Cx8m?%x��6z�r3�
u;� ����%yPLi�����3`�Ʊ���P����L8}ԯ��:k4R�3� �9HT$�v\G��@��,��MD���p�D��Ȩ,��o�$�/��(��a	��z>"��R�ʭ�ܔ��Kaço��~��2Z�j:����0�z(0	�4T0,ӻ-C�Q�Bdۋ��K.�ڿ,�z��﷮��\@t��gt�9� �a"�L�_����}sYI8��t@��f��SR�?;j���4{�dwާ�XnQx'����\����=��_N�L֢���z�Y��3ٰ��ÿ�r��V���c��_�`�77��ew!giCn�C�S8Y�>/����@�5��Y~����!�����`�F'���!�Bofک�K\?�K#9�Ӡq�պAו�ēΕeq�dSap�x4��T�]�����P���EjQվOL��X���������~�GU=�O��Ȩ�A�ѧP�\�,�j��c����ih�;^��� ɾ�����*�D����m�}����(⮸�!��ܵXS��R\���Ib�U���{�R�	�W�nn��GK�B�z���[]��������Q�f���TDd�6(XS�u� ��^�u�}<14�g��'X}����>�/ߓ��'^�ĽI�)�w?�8��g\��.H<�a_�Y���&K��~�1ғXy�kl]���6��՝�`]��?S~��� e�+��^v9�d.
��*u���eȳN~S��A:��"��/�&%i�Jb�f'V�;Y����f�k�u�v�� BяH9%���9'tn�\�ր��we��6Cv�G��OF�����ֺ/���&iA�(Qi�0��N�
�Jic�/z�g�z=��y�B�G�R-||�r�59���ԑ��N��~ډը�94L�k�
�k!�o�5V8E������oNN]�Uwp�'�-Y�J�H���;^��ި47_�[	���U�_��N|����Nˢ&�%>��b�e�vڌ�^���'��p��V$5�P����Em���^6�5gY�>����x�)d�2sq�}�F�B�?���#r_)o�֣��@n>������f^��֏܆�Ȇu1��s�F\b����V*�P`���^
�9�.�2�FG쥂n�`�#u�Û�w��5��a��������Gs�O�w�ڐs��i���[#���kd��fm��LZ���*^����&�v.���A%q�6�!����hi�� G�.��|�޾�r�R:����٠N����lƨ����o�ުaBS�J`
���YLK�ܴ��U���vƋz�I���f۱)�z�������p����Y�ܣlX��{;��ge�v�bN,V=>/��ty
"�!4r��[�W��z�.y���u�?{˳K�&8(5��ǲ턕��[�߄י ���]~�X�<�p�#��*=��d��N�����H�:F��s0ݻ�`���U����q~�J/�( [���Ar�s��15׍=_� a �e#s�7�$���b��<А;c�F�9:�w��2�%Y��zL5o�ST%Ѩ�A��F:Y���==����!����S��l��R��M���yy��U�5~��mMp���%�v0��sݗ������R�/&CP7�!ؕzhQQ��^YYbkJl�j�<�����y��E��
��LI�&x�8?�*��؈��]�G��	���19� ���W�[�2v%Z�+��WU�a2dĚ
@�̅��� ;��˯(Y�b�F-*�ޜQ�W�!�uҬ
���mWPP����)�aoي��q���)�Oj�pc��$�N���ʞ�3�i\�Y��ڰ#@���\�g����:��*&���N
=v����/:M7�k^+�'���U�f������iZͱI&��i/N_�<Lڶ��]�j��e�>joEJ*���o(���=h%嵹�E&�H��I�TK���qn�IJ\I?��%�)��ق�?�&ם�$����1��=��2h�g������b�����\(����P&)1�u��:W=RKى}��Fԣ9��y�ޱ����i��3i֕N�ͭ������純�r�.�`$b\F�Į��~QBWG�A��e��h���ȿ	��ѹ���h-�,5t<O�k����X`�n�b�>����Y�"��"��pښ����0���'o#�N��"�v�G��u����h�.e�)n�uՙ�_T�"B1�J� ��xI6f�?l�����7��'��[DH���.L� �G�=��*=P��:<��V2�����TH��<蕹τ����|^�y&�x�4!f\��c�C��3�g1~!o0����8��9�k�`2"�";�H�&"�>��u�Z�꧟zq����J�̓"�m��}�`�t��e��+�9�v�A6�����LC��ZK;�Jɮ�����S��TZ�N�������E}��{x�()���*�:_��Q�RK��k��AT�Ē;������.[M$-�������S��K��îu`;TI�C�ƅ��J��2 3���v��0Kg�ԫZ
_��%{���A��]�&EX#I^�%���i���~?��Md�� ���<,�d�t;g@����z/1I�ڦ�4k�K-:& �L-�x�)m��n��4\��Wjꮥ�j��D�@��w�`����!�َ 7��1�k�j��lya�(�M�e{���(� ��K�Ӵ^�wb�鱉��7��-�|�_���~�����qcF�X�c���� 3E&:��T��FV�2������
�q���1L��"���2�.\OǱu��r{����b�����TSya�DM�J�?�mM�ԃ��Ov3W��{Y��3�V��h lƚR!V��l�6���&L'��LAf��L("��p��k�6r�������C����P���>�'��e���pp�Um�u��?��y�ѳx�gV�@/?����|�)ٲ��|���4�l3g�~����c
%Fؽʣ�";���W��	�O����X�x��F��n���N?+w0��������FA.�]]��T���@@�� S0���u�-�PݹXof�����|TW�oLh���YT�j�Ų
�qr����ߋ�8\�"�����.�}"���PGqٻ���oT[3���d�e���!�s���fyjjm{~�y��]9Oz�Jē����>����	n�ΧB'W����[N�x5z6@Q��E��C��M"Au��rX��j�\9��&��d�Z�pmgĤOE2G?U���(�
_��>JUOIO��ni�s%��Շ�z̻=�4�2|x�2�F1�i��l�G�Wc���7T �.�Є]D��'�gʼ�/�4�AR���19����@i��&��_�:7&�;���^䯒zm�+����\�Z��6���ɜY)<uL>4����~kY�E4;φ�Z%����.!:��#/��*Ma�IQ@���dTDHH1�9Nch���W޶���;b�y��38!h��	c7帓��|{w����[��g)c�b�_��>BF���<u�����=�x��(��;>)�	�<g����D�o	<~Bl�����ҷ��h�m��U:��]���V>ȸ�\<��qSm�WXM(�+�DOd��P���	ezU�0��c�7��1x1�>	������9q��@<C�����=������p5�yV���P%HZ�OϙT��� p���q���E�yЬ� �ԋ;�P�*z`K̹�Bo�i�i7�f=~��P)���-�3�`[51�k�WF1�Y�Z�DO�2����)&q%��1{�"��E��.&��ǎ�Xry��#Iu.��zs
t�I��EAۍt1�N��r�{F�Ǧ��O*9�6�ץ���xnm�'T鬮(`��Z��D�&{b=�;�7*�b�^����f��P��i�ҋ�����O�Kp9~7E�n�!H��P�R�#��QR�r�ųܹ�^��3Z�I�����	��ﲠ�:��x��ӕ:�U���c�p�}dG����c�x�g��
�é�U�	��	��ǩ�}V��T�O�8�T�s�l*�9� �gF��Gof��b�4E5�(y�G��qGFaqa[���Y<>HW�:�NfS펄�S!�����Ѻ��,��ސ�7��~}g�&
�R��B5�D<	Z���gB��ɗX'����6q8V���6�C��aF����i
	q���q)�hF��ؤ'0��F�*�}�]0W�F���S���O��2CQ��6sF�C��ⴝ�G���V�'��m��|}��u��p�!L��r�k���O)����2rI@bXUӌ����;�$D��8�W�t�_f9o��֖&G�e��NUL�p�e��T��Z$���a� ��@��^���>j2%�v���'�X�o�~���3l}
QV�5�]�f����s�H,�`��TZCZ) \&5�!oޙ��+��d�G���v6�%m��sq��]�J<�im*���Æ��'������Ʉꢙ"z�7�1I,�r�� �=�Ԃ�㭀O���i^
d�X��)�.+5M���,�A�1=��{��Q�X�����jj4Ѿ�X����5�l^��Ô����A�*�{rfS,�,��6@O8���ğAӬ��� ���N��dr(ݹZ�d��b�Trtӎ�e�}�6�Ui�c5��Ei�93�
ۊh,��lc����pgՓü�]��%��'��L���&��?ar�mbv�{���M�)p��@qLXA�T.��:��׮o)�wPD);�R���'@�!ھ��c��g.a�o��JVj�vZߌp��_A�)�U:tA46g^�N-��7$����R�
�5l�6�]M����B��^0��5K�'*W��bb]��YhEG�N{Y
�B�J�ͮ�]=n�j/݈����2f���@2�54j!J�[��d�><�0#�3��r"'=�B�4u�&ۇvT���: �L2m�K�uZ�ν������G�t(��6�<a�_�2�Fc%h��A�	k�E���'�O{S��4�՟�ҕF���v�+�j�l��i+���5[K{���i�y�c�� p�j�FqZ��/F\E���л��߳���H�m�y������<�F��g��˼C5X`˝Q0�<x�_� J��o�L�F���^�������;��ǁ�ޅ��j�}��9�FW	1=�nP�p�x'fj�?#9%E��K�bcf)����=ʇ�Zf����g�T�F~ZQF�6ۙ<u8��4?#����}��F��Y	z�Y��; k+�@0"���Ne������ƻJ���g/I��Ɏ��+$�y�N�ʖB��|A�Q�r���K���������l�HGy���A�;����N��;��hT0C�US.��"�A��[v~����~��o̦�tK����ȯT�!z����N
/����O������7&�q��4_Q�D�HN�灾k-��h�:��p���m��8*��ء+
�#��E�t�[u��Ü�<��ەa�\������؞�'2㳕H?@4kz(9����-�����W�+�� 8ܹ�r��o�J�m0�g9n�P�g#�K웿bPM?u͏���~�"A� � ���33�H��fq^㎃WvZ �\+��0+�DT�/�/X��u�����r�\[�������uU%v�͗��̀Y�yv]���a��q�A#�9h:���;Q��dO�/@���\]�<���Cs������Z��ɫY��ԷtS�ݫ�D�(�o�Za�}+�q�KE���ryeX�x�&r8mp[5�����}�Ph��GC���9�y�ըtʨ�b.�~������D�J��8YE�s�=⎺�ߋ�s�ږ��Z�eIf���.�����)���1�N�D셧1�����P͟&������b��23�QQ��O����si�֐d:��W ��ײ���R�T�\s����K$�q@|��W�S�	fa.���z��hU�ו��5�7!<��k+���%�@���B��ļLrL����T��]�K����8̶�.=��SB��պc��;G}�]�Kg����-�c+@�qc��c�?�.����s�+�٫V/T�h�/�7c��yx���S����4�<�s�t20�л48N��5�P݂���b��S��d���+k�(.�S���Y?WjTSc�t��A7��Cږ�UT7�)�<mW��\f��jA��n
D�]�Ie�2�jܩ1�"�`�vl-��]�[�_�[���Z�1��m���M��ؒ��� �0��	��&�(R��kp}``�_a�k�A��s�����L��%Z�+�jeח]k ��q���.�j2����*����F�_����x����:�B/��t僙(˅]n���TmJ K	Y�#��_d�OU�W?��I����Jr�����)���8�M̾��l��E֧;d+�A�����\�|��Ax�H��ʐ���ig�W?2%���� �Ƃ���Yx-�I.�\��6Tufb5�X�R;����rW����8N��w8��[e!B�b�!V4�"?��u�£���_��_��G��/B�0�#-���2@�0�E�����4ˉ�d�w�ӻ�/)TS�;�'��mV,�'����	
سe��?a;�hL5�F�`��f�&]��)#�]�'jC��?[:������ųV���X|D������?��R�9�Bd�Ġ�t��h�y�~���	�#�vPpfc
�i�t�8Z�a`�P24R���9�e|��Ka#�#+hv7%�	���{U9�g�{��Xn2�~�0�$�\�8"e?�֬*k��v��KU�1m��OJ����[J���ǿP��E�'e-.�;h�9����;:�3���;M1�Y��������6}�DAڮ��.��U�lS������T�L5U[*f���k�=���I�{�|Eh�1����'�O׆?x	�ސ_���/,���y�¾��Ff����r�LQ��CQM� �8�Ӳ�d7y��<����@߮H�`���8�|7�P"�O_��,�/��C�J22��z,�:�E��*�F
��(m��I'qJG���׷M0=���RnN�@/����-��󨽥��/g6����wL-@�%�]���A.��~%�f�@X8�,�S\I�%�spZ����4׭)hS�T�E+vq(�T�	�?S3�(`����]ə��)K�]��`&:�~:���>��yq4���H�m���~'���Mp2�mz���7�)���K���o��"�}<�-�*|�Ib�|�EL��c�b��PA��>P¨����8��	��.��]!w��[ M_������0�Zi��B���E�x��h��z��_��Տ7�md a���S���ulQk��[~p�A��o��]��	�n��L��5��/�ꜟ�'7S�1� �������l��ŹU�-7o�t�ܸ�<䝞��4�J�7S�8.�����j�0���[�f:d���}A�����@<zl�u�k����!�,��"4x~�߫דg{�_ON���֯
��������bV{���`<^M7�g
��g}\@�'NE֫�v�)�d������O��#	Fv�؈�8�c!k��S����[a7F9���w�&֛�����6/J�٠�̈́�iS����-�
aVgpH=���/r�b�Qf�x��x�F�t�"¢���Db�`h���
�r	����M{�=��=�t1 EWe��P�P:��D�4�ã�'K�����]MJ.X�O�M�g�+�S�
ajU �w�=$}�#Gr�!5d��ē%�~�Z�J�JZ�ݏ9�}���-���&K(�K�k�)//�bZ���:��i 4��kM��coKa��p���\�nDM��#�A_��$�Ģ��>��t���<�he�츺��-�tVW�����lm� �GW+uG������4X�zo^+ZZ��j}f�3�.�t%=�G�\������A��QW�G�c�T�:�[~�6|�A�a����[�#f����4��WJ5�p-5��=e������IA=�2S���i}`
��;3��!��IK#�.Zm��ġq��S�m��2�1���^�U{��ʒ1]ʺ�*cu��q�0RZ����ފ�r�Z��"�S�G�3�$6�p�42Qفn�b�ԣ_�C=�!y�m�|���,�IU��a~dp�};�2 1�/ģ�h�⢮�AE=�$�q������ ׿�¾�j��V��wW���W���Sfd
�����.��<��
��0ՙ�}3��Q�)���Anc�rO�IA;���?$�)RӀ��Q�a�<,+�1�dL�tTP��	+����9�J��߭�ΣD���	��ER��b��C�����T�F#Sމ��	�o��V�G7bj����q�
<�Iid�"ڟ1��US!�F�<1$Q�+�D�`3��\Q,9����"Pt���d����\P-�*�Ҝ�0
��l��Ϯ���SU�ovQ�������׷�Qj�b*g8���}�c��:�i�?4l9��(�R$��'�7I�0l����Q鲙-�(7���.u�ܙ�!�_���ڈ*d���]�G�|����֪�C�ݧ�5��kqi���ˡ���@'i����uR����HOK7�0��'.TV���YTVFЕH{.'���z=��:�R-^R��(�g\h��n�.p9�c����I�3.�:����B���]�=2��^��}���l��oN�03�닻�kG�Bտs�%�*�#Î�{z�F� �j_�
"�[<Q1�;�d*�^ B��ed�V3r�9�r���5��ǅ�8-�]�D-[f�	,zW���C�����#�1����܍�Ǵk��5���&���ڷ?�u_����7�R�
��ilU��wW�5�1JQ��h��:��Ua�m,���y�55�mK7%:(�b2 u��!H�YX,RZ�k���:)S|��l�������z��o�����Q�n1�T���q2:]��(�"灻�N�Z�r�]��9�˄�����(���jT�IP�)3b���l9%�#�~k�
������|9�����/�u��9^�{�p�N��� 2V�������3��"jP�\�p����������($�G1�\����� �"�����0��'{�����O�-������)�7�|b����a1��I�W�1�^��������׭��:?��5)�g/�?���,�r�|��*�O��NU.T����)��íP������5m�j�I��c(PS�`�Ǯ;����D�X�A?���Y��KᏬ��>��A%�]��U=\�Oi6=(�?Do�fWO�w�+˗�r����J�Y�N���7UZ��ĮE��g��E]ݏʱ#���چ����I��닖�*c���z�R�ԑ�˴���N��x��JW�Ц ?�t-���w݈��o�pL���mpȍkJ�(k�<>i!Y����m�=|�
v�+ќ'��Q�HP\���'�ő��h��wN�!� 6]�ZӰIϏ�:��t#�ɮN�س^c�%-@��q�jxK�%�$��,M���_WSf�H}x�+~N�2���%^|J2�y*B_�(����j[`V�/��:�M�h���Z-b�``�Qs�y��|��݅��Bo1#:�?r`��X�?�aK�;Qo%�9���$�LCO�k,[�\�n!��=�tS��G�`��'y�a{Bh�����lGm_�D�./�R���2�W�EU"�{��v
<_?��kk�Yf�ʯ�i���%�2y.C�/8q{���̓?��t��q{:;t��$�T�	��\B=^�auR��39�x���heq�Ʀ- ɸ`��R�۝���d��y�cxs��jENV�e/0)�ٶUbT�[� �
�h��jZb�cy���;�\���Y�u��k�oi��+վJ֬�8�Mڍ�0��;F��/�^��2�VB����sO[�!.b����@g�$2�؝@�]�O����t�I:���d�>�*r�X .q��P�_<�J
�7s?�mB�Pۣ{׌�I��O����;���a�^�J�1�޵�N,��M¨V�{��QΟ4͜"'�anO������ ����|hoT����xR��ǎ�8���'a��6�7�1��fj.,3��.�����n�7���`�9.�d�"/^\[����&��Yo|��=��Q��l�çs�ߥ�I�4g�|�	�7P1_��:�����Ф�Ə��"�W8�ll��pk<k�	�+����!x6���L��������{6�S�!�vt��[��5n�U�� ��<Ĕ'4"�^����xsu��a��1ߊQ}�+�J?���Hwf6E$�7��C��[�zitj��"�-��ں�ˠ�z�l/l�7��}!2��Q\v��5�_%g���8�!�yIe�X���^��"���C޻B+Y�.�z��fJ�����9��2��Z�u\��@g_�?���GT��oZ%��,�ىt�_��5�gp��%�Ƙ�!3���D����.���;�b��⸼J�b�sz
6{�r�� ���Uꞣ���R�4�K�D����ّ��r@ ���9b��2�����0ng�V��ջ��-|�f�+P��R�>�����M5�sN��H���6d�;��Z�R�Y9'�R5�
�]~<�������T�Hk�+6!��Sn`��I�~���e4Ok����$e��U�]毭��m4?D�� ��U�������7����ٴ��m�\��t+�Wt�7�Zv��}	�!�
~���tZ[\P׫dм>����N�����'=����H4{�a�!�7�8,ە��ox��f��\%a%S���L� ��-���ê6@��3�a(m^��l���������U����W��j$���1�����(A��vI>�O��}����f��Oػ�T�|��V��)g�20��_Q9�q��uB�k۶�JY�?H��+u��	c'w:;����Rݟr��2�m^�Ϩ�:r귮��փϜ>���@7|*O�F�a&�(��U(P�	FO���)�����!���ՀẂ��@�d��S�6s'}���!t׃���3[�x���gs��Fi��=����"3D�s����T�Yiڙ�w�z����z1�&'�SL�5:�o�z�U8<R�KH��Q+���k� �"N��#X|��S�` |D�����Ǭv'� �!�\#�ȠZ�.)�/:�ӖC��v�N��&��d��E_�.U*�<GX>��&�缩rF��ԗv���r\]h�h�-��L/s_��#0ի|��z��EXd�e�Z�=�g����B[������ �d^΢'M4i|�����pP�91��x�³<'?�ZQ��j������sG�đ&J*N�p�X�;�ty����d��y*|�9��>�,�t��j�-j�X�Y4)��^�RPC8�����A*]F6p=F�"Y�#�7z�a��	��>ld0*y*���*e_� أF%�y�ڟk�tS�xAe�R�Z��?�=�V�$�J�q���Q���z�!v4 ��C:�͚��>(�7�k�E �Ke��m��n��Y&`���l����E���*5
~��|�T���l6b��'���G�.in���\>J���rE]Q!"���V�KC���M�l��Q�e����D�7��р9������!�klV�����la���"���[.�Bb�����Ȝ�~�ʆ2j{��J�#��5'�ؐdk��\��V��6�S~Fm��,�>t�
��c��(YUSey+�����^ I��!U�sm��[NW���=^1��=�s��ڳT��u�����d¨�ʑ5� ��m02��K��~��q���7b������P��6��	��R��γ'9OWob|��R�_��J`)��!��y�@��������N����@a��*�z[�9�	C9�i%,�_5wv�9��*v_sW�`ݢTc�|�?C�ސ���tz�-�&�EA����#9CXoY ��Ϝ�%r�=Y�,��
�V��]�c�5����HЂ(Ci(��0o�|5q�����^�C�0ѷ�?01V�Gle�CFg(ZF2�/r/�9&����b�Ĭ�B�K�
��9�o���y�r
W�]��5��Ba�+6wr|�D<�QC�*����A��e��F-�8�](��*��b/ف;�W��]�G�Lm�XdZ���^�W江w8������S+bdI�]����ħ�L
gC/�Jzw�7��A�����iĊzoy�0}W�*ҰE�$J�(MԺ"��,YG4�>�Q����� �GXYeS��X�K�t�U�;M�o}���y���Uޜ]|���,U+ؚ�#ë*�!�|c
�!������+oy:�51��>A����gh��zLL��5Lh���U͉��o��~���p����M���ݟ����m6{ׅ�:V�:)�A�q°Eek�(i��)�B�]z���:��Rl<�dE�Z��F��ײF��N-Ig��^�� 4�y���8��C��_}��Y
�D����_�5	$�Z�h�1�+`�)}�\�%d��]}���&��2��E��)]Ѳ VvJSEn���`�d��H�'͘m����o�٥�s��t���ge�}��X,<���[����f��;�g`���[eRe�D��Z��Z���d��;����(D�����wڒɛ+s�f�z�~t�7���;Q�D��e)�s�w�s��Y�Cp��1q}�V��@/6��m�Nr���𐔵Ly���(���[;�+���9�������o���gX��[��FH���	}�����`b�jK��/�O�͛w�� �gN7��Hfh��|[F���w&#��	�)��!�:�.\�T�B�MX��:F���Ș)K��0mqt��+��F�_e_{1[��0NXç��}��"�?��� ��Qa����W�����v�c
Z2����A��-�.���,��\�+��+��m�^��w�P��^f�F�lи.&U����o,��#`-6g��d�����2�J�W&2�*��<�ʚ��`=5=|�a�E*�F?<�ⅽCo�n�^�����ދ4Ǿ0̸@@��s��a��F�[au�֤Jj�q������{����%>�5���_XH��L��*ԙt������ZDd){��[��L%�\���-��i�����f�YQ���Iy֓qg�/��׸\h���$�ȕ��&G�@�0.L��Y=��K���3��;K���\�ۗ�J��g�)�a8�ߤ�"+w����5'Y\O����{)���`6$���$!�+����������q��w����Go���4EK�*w�[��:sg�;�z:�im�,
&�Ov�ܣ�I�ͣ>����`�z�Ԥu����NN٬�Zq`4�55��i����Ұxa���?JT?d=�x��7��k���6g���r'���)O�hW/O�����ܵ8d��X
�ef��=+6����56p� ����YA���F�~���6����D/���������Bml���s��ɶ���#�W|�����̎�8O��3��l���n���ư�E8̞R��3�
% )[�. ����d��'�C&t��^��Ӊ��ؼ���XfZ0+�Y�hq��D��k:�V��s��6M�{�����X~��9�b���t��Я"%v6�A����$ݢCi��d�_B�2���췏1��xqs��Rs^K�����0�0iHJq�c�d�G6�W�o���){��=׋ꦝ�
{Z�%������V�E�Z�4)�_�:��*iI�Gk�R����M��*��|������/�T��՛��;����J]��=��`�?� ��3��yH0p�������_�.%�����9��Ls�&2�8�Y���M��j�9ᾮ]�)-Q�v\�H-�ME\�)��Π�ybֲ�7��Yr�X�5L��s��g ��V��e����v
��a�#��Qɶ��`ͨ�פ¸���s`��#(��V��� SH�ݒS��a�b|telPdc��_x���0&߮�*�`|��5IU]6{F6�#tJ��j�h��3UĎ�*�f��W�
�8�����k�a]�Y�Xȧ �Bq��z��$�]
،�M�/�k��Lc��� ���l!�G<#���@y��������w�+�?��v���t��
������C��~5H=��kY���[ε	�����"R(��0s�:+9�$�b���D�3�ڸM4ϴp��3/�&Џ���\y�'��mӜɯ؞��]G�`�ӊB:y7Q�Z�遄�;^!����*��#��	|<�{���Gqy����m��[�\JE���+ڄ�_��B5{LXI:Xj�K��`�����6Ho�]�Px��,�N� �O:�s[�i����'�n$AR_��]��N��?T��os�v��z�Ӯ~o؎�'{�c8*V+�8�����m0"�8�c�3������{�aCU�{���I�=�л�@��k�Ee�-a�s�.���W	�Bk�y !̽�G�+. g������7q�6+���T�=�,��Ex�N�қ=^�HMKAzX�&�4��F���4��R�˯	#-~U,�A�A�=l���ˣh�ZUc��:��#p] ��_,�	����Mq�~�F�ڰ+e��[%_� 8J��z�h>`w�!܌�Z,4n*|��J	pZ�(O �e;�Tڤ9���	�5�6?_�4�3=J@��!T��j��N��m�e���}R�����芦އM�]׻���V=@I��N�#�G��}G���f�^�eK`9�Z��EϽ��TI�CsE`���g�8�mf��ܾ\��@���Eգɦ-`O�r���`�NІ�gR'�!Ԓo�Q�:σ)c~��ȬL��(��M`�=_>�Vv�7�p�&��O��X�JX����L��0�p}ŉܷ�������uU s.���˫�#� �C+��/����Ύ#e�{k�m�8���M��^yX�1�%�V��b�#T�۬�P]�������7���=�L�\?�Wk,Zٸa[W����&��gp�w`��o���(:_�զ O���>��g҃@ױ��9M$S����\�]�{�Y�\xKt�]U?���u� Ph����K�R����c����j�$Z�ǵ��$��T,p��/�)EOs��+}�����z==$���6�0l5�P���g�7Ο�Oq��z|2��$U�D٦e�����
cl4���6S�f,��P�S/�k1+�y"����\�k#��͠t��`r���.��~��^9�hp�Ȃ��6X�����U˞W������h���
��=���m\f�L2(�4��	p)[l�4ݟB]@�Bm+c�.���Ӣ�6�ꇿ_���lA��me슃O���ٞq�����y����ꍸ�CK�	n[�0�|H������L:B���H�����
KJO�+q�SJ�3<��8���	�����fE{��0l��o�xO}/�U����A[�:M;��^ķ=�+b��)��	ݘ��'��p����..v��1F��c��_zQBW�Ӻ�� `篭�˸$��?�8Ⱦ�ʋ���>�i���ʿ�"�6�x�6���-ȪK���,��=�{[�N^�wc�W�xa=.��Os�sv���V~8=Dިx�o.pe*߻����= �:'�Xj����Ṁni-��Гk~��*pΰu���}y1�{Lؕ&��1$"�R�7ܔK�)��P�ʤԗ���[��kV��:��Cʑ��i���\W����$�^?�E� ��(�)h.eA!���Eu��m� �BCau:u4?b+�����n� �)Y�VE�	,φ[ag=�>��㰴����nP�U3D_w^Oy�X���`Z&#��ЎP/���h~��'�%o��3��x�q�9���xP~'��8Ǭ-|
��ݩ�|/Ti���^v/L�eB�A�C�7(�i|z�~V�d��^���8#��Rke#J�.��
��vĀ����YjM�݃I��Dg���>;���I��I7T(-1Գ�&��l�&�rߍ��=#��^��+>��k����<�4�q�D_$�AA��P��9œ�Ǉ%i+��Z��!����Η�� �[���?����|:g�	)��(Kl��@�uK!-�`�=�C$"�Vt�f��:�I���/�dZ��ԩ�ݾ�`
�u�Bv:?��1܆�n�Ө�&�
xD������_�Xa�[t�ݽYQ��F�c`��Yn�/2 �c]�#Wo��,�n  �+��
^nL������0��n�겗l�Ō�d��1�hy�
Cͥ�2��N�h�C"�ˠG:�{~�ȝ�$<: �t�Q $���;��j;���d�Mr1�3�I��=�B�d�Wa�3�sp��� -؝Y3:�A:�)Qn;��2�_'*cJ�]�i�lC�Y��E��m`Ч{n��L�+_x�P�!����>�?k���Jg����|_0ɢJJ���7�s=�G��#��Gn��^ J)8H5+��(,Fw�Wqcg�Yz�'���0�S���ŏ@G�ާm��D3�| Ӧ�\#ø~��	���˫-����00<�&4�h%7,��Ob^�Ol]���K�^�ؖ������&@�'�7�7�O��h�������S5ѫ�&����f�ΐ[�:#�=��I�8v���= ��nX�0��O?4�s	^�&�G����R�ˬ]=�Ri�(�+a,��P �:��'��ј>Z��zqA���@�<U����'���n�5��#�6�@9I��JJ���oPҍ�>)���@A@C���V�.�G��q�C��%�z<0Qⲹ+�|�Z$���b��?�n���ʜ�vg��=dh����1m�b�M��U���0�ޒ��M��4޹�������]UՋ�zrI_#���%�Bx�+�,z��/!��%;._v�ǣ�9�?f[j"�E�ʻ`��J}�<��!*l ���˜N�)��^��g�� >�������1����Ɋ�"����(�g2
w��W6Fd1�v���F^�����
��^yѪ���fǀ\��Z�����g1[ct&ې�����"n\��\���i��#N\��+�_I
�@݁�O���3
R좐�0�O����^nf�c�������x�s���c�#�Z�Ո}�H��m��<�p7��[`%�q�.�^�@�͎���.�c�6#_/\�ڈ��i����q�/�H��ɔg��z�$Sm�m��#�e�ɖԭ/Ƶ��v�"xY�WM`�� r�Ź,\�h}.�=	�Ql�Nye�����^���D>�3y�l �:�Q�����@M����ǎZhN��Zf�1�S+{�8��-�h�D���JS؉�}Z�ʩ�J��nt�ڵ�V|����ZCU��4+{I�������tF�a�<�K%��x�z
��9�k'��v�'U���[��@G�~݄����=�8W�^1�8�{IT5��&�pi�=�O�#�4I8Q��ȱ;�<D�t��a�tX�W�]�l�Ky<55Y��|����.����W9�{
tc]>�/Y���lCJZ҉���g%�����|��oi� �� �ٿ���T�ް���U�E���B�
i���0�J�<0�j,����������f�==��0 �4�m*��c���d%�m��/_�՘|�����2�зS�Z�<ݓg��=j��Fw�̐���ɟ9��{�w����|1�K�T,�U���E���x�2O�	�����dck�������mm�ⵋ�tL��#|(��R��cU�[���i�NW�a6��lK �=EO�Hom�w���<^���W�Ǵ�2���(N�-Ъ�/�jgW�@eg���$B�1�"!��?@0�KD��d�����v�hM�pe��\ϼ��W�������5��˶�w� T���:f��S�Q^��@'�޸-A�wVg��E�~�h(�e���|��Z4{�A�zB�s��M�ձ?�X?�s1�Ć�HwÞ�[��3g�\<dQ�'�5���/�!� �y��9R�S����GdZ�nj]��~�i90�3Ye|ϵ���XB�b�.N*Z7lOڷN�	D����aҰQ>l�� ������1O{����X����R. ko�r܆�U�1QW8{�c^����8�aXT�P��F�3��� ]�G��+��"6HDZ�Ia�l m5�&Un����.OOE�����6dϒ6��1�>MZ��|R���?Z(�ux_�G
���Mr�u&��59��Xt���,��|W��ے�4�n�^�}��d-a���ޙ��E����f�M��r��Р@��C�{N�ƘP�h��NI�j����\9> 2D�U���\����ϣ��|�^��L��Uk�E�ݺ���j�l��+p˺�a�G/vt~�Ϲ��؅��K� ��>FrɈ\4�>����#6һV@�J�
�:������|dv���,�p�!P���m��f�Cw����6���2A��L۵�ƃ��Lg�c��~�Q�2ER�@1�r�<��~`�S馧G$'���A:�F>����% ���sL�o��o*.9���^S�ac>�^��p��ȅ�enw�N�c^Ɋ�y5�'��D�U �Ax6;�bkk��V����wI��t����G;��6������y{�*b`.�����۽�N�et)�~�t�{:=�ZN�D���Ǝ��5m�6t��xwYi�5WR�B�"O�iF�v୙��_m�&�3�U��i�g<�GO��-���;��0���V�)�~al�0zV��Z���4�R,Bn-@P�O}c�Y.�/ >L ��`��&w_���)�qMd�'��л�J�)[/����B5��4`cM�h�����y�$0wL+���$���T���D]W����M��EqM�,�\�;Ti�p�6�
d>*�.#*����Ԟ�1E�jG&(���R���.r��2��ɬ���S�A���hӬa�8��f�10�G�'��e������m�J@���/��q*��V��BH��R��}��J@�Q�h\]�[��}�5?=m���E
�9h����.s4����[Dm��[�m4�r��+ڦ}B��rӺ�u�q��~�<���X��HŪ����C������œ�+%잕j����C�y�q7�}�y�粕���� �!_x��������*�����X���<-��1��;GiMw2N0hW9�]�R��n����S��#��c#,Pr�'���cm�",T� ��o�,�4&-M��m`���S�����=pz����Z()�pӳx%��+����S����Fݕ���-2^f��ړ�c9�pu�$1����?$8��l�orO��m�6<�6+Z��r�W��;I_0�V�-�H�&Z�g>��R�V���Ǚ4nG1��w��N��mZf�Ԧ�����qH�>�p[�Bp��.�b��� ��M�F�zmr�+��\�<r䷬�A6`���໓��+��Ƣ��-&$�\e�q�rc���Ɓѥ��_c���2!�`[I.���T4���� ��+�=i�M�^(xF�Q�9�C���O�4В�'�8t�4��-Ђ`�jm_�g�a���n-�6�}&��WP)�*7sm�y±�G!��dAN1|ƭ�c��Lb�NB�v�%�wY�Й}�h�Ƿ	m��uM���y��ٸb�i>�Gf���b.Є��3rD�OH���������B�٢7�铈���E?$?`H�_��1W0�E]��bVw+y�o2�	�\��:
�b�<���v�O0!�)��@�?��L��fɲZ�qӯ�%��j���GNg&	����k3%Y�@4)QpI !@|�Х��]��h�H�Q^�E$�%�R��9���ٙ�f��x�^>p�~W�Raf�y�l�E[Ye[����m�S
9�	lx�����TG}���&L�2pj5�]ј2#rp����Z��觬������xYݷ�k^s����k�L�}�8[��/K���9�6 Fl�Ü��}¾�"���b�4�C4�{z�($5X��2b2bX��o����M�1x�Dw'I��J��f6^\���Zd�Ѣ��G��b0^uY��)��#�l�a�ɹ�_��%��琯���z��*D����l���^/MA�)�fr±��>��6�!߄�v�&^F�4�.�Zʰ�Ɏ�qq�q���i�'8�*bT�&(>ɝ���č�Z%k�mZ1�B(�D�ޯQ���N�#�f�ȕ���l�F�!����ff��}ܘN�Ђ�K�©�؋����Q�|j��@(�ç"�1۾��[�~��B o��;uX\X��>�~�u��0�c�[�����'�Lc6uJv�4�����ca\��Nzش�����	��g+�� o�Z{����:0���j6�ކ O���j�GFuL��a$���|���W���;J΃������r�ZB)�詗�D����C<�}ӷ��&���-gy�j��$AK�n�͎�r4-�3�O��%;������x���[�����Z�t�l7���A3]5³��[m���8��Ben�*yd;,���+}7
8HjbꦰIB��&�m"k��<�r}Dp��P�����E���3 $��FTΒI���rj�g�G%�ک}�m&���[n�:��@�͝屃�s�95��@ڳI��a{��8��)(�\�(�0�����]_��U�\�m]/rY&�\���%H�0	q^{oO���iW��$T��W�=$��ð����o�(��Čz�k�T��2F��Jw��n^7	
����LI�J�C�*����@Kb�W�h�-6Ϛ=���Ɔ��
���Ag7�t��@�;���u2���	�����Q�P�j�C:��O�q��\�d�IP��܃�"�� ��v�(ɍ��s�}c�Տ��QK��-���F'�ﱯ���^�XU�/��Q�e�n��ǆ`̡�?���A�o�h���)��!�S���D�W�T���8h�߄Y8訝�Tz��n3ꮒ��@�_X����h=���8��{�rQ����s��6��ʳk)b+Z���9�$�Ihl���wp9~
�&��؝��-29������2C��y���8(.y2�r=�wy��ko����M����E�#��1�����(�3"=�Bk��5xd� �X����ط����v�ٙ�-���`�tL����Jm�w��[�z$�j+2�#<�/G�c�	��յ�Ϫ��A��Փ0,\uj F|�o!aR��s����;�����O.����mk�;݊�9���N��U]^+A��>��)����#��q��JSY*��ɚ�5�7t<����rϭ��{#L��yxa��Bw�\�J�Ρ��$L����q��*��S]T�_�y�t2�n�ڠ��Hu;�R�tw��X�Dr�C�z)�kf�8�d��"���|����b�j�?�!힚{�|K����Js����6�%+�TU��C��>�C����t���*�U�}x\�N7�s�s��S�?x�.���|���Q��;O�:�~R��|a���`��
@2e��q2q�Q����7/����
�83��{̕�x�����R���ꜵ]�ps�|A���|����8�Ƅ[Ç ����B�Շ����Ta��p:����nJ�Cm���{�O�FDs��ȹ!ո!�LE�������Z_Ѱ�9�O�Qa��M�u��#��`�p��u 9�wo�tC�x��&��y�>Y ����5N��i�@�$G�`�Y!O	��w�4̪�Tq:E|�Y�+c0���y[n��S�v��2�u�'���pϪ�ɫ �;�'b�S7�N�rQW�V�9`��<m%�;��
�:�"�NFs 0�m��^�7�Ƃ�
BH��z�%q����G�a�cPл�������S��p��?<�S�x�BPb&�.�tc�y�� ��~�Qi����G�������	��|�!8ⅷ%�.Ȓ@S�%��,D�G���-�~]?B����L�E&�Fnn��]O��'�tGpv7�?����Y������Z�\k�R�ѧ�2��Q|���6}�/�"�/O�+��4�tv�U��%*.�u�"0B���ުmy ؝��0�CKV��C�p�E��|¸�I<|.�{���I������9�c�6d�K���>�����(UQ���?{0o�W<��� sA1�o"�a���)[�щ��Ɔ�H� 8s���׃�8���Ro!�/���f1x�c����H�ˉp(�sJ���@x<w�52C�b�
�u�'��B-�/��zw�C��L,m�TGms���5�E��s�
k���įx!gA~� �r-�p�l�6�\짽�^,�P�➡z��rePT�C�b�Y��B0���<�eN;`���B(-_����=F�-��4\��#�s�
cq��M�j�Q^��m)�9�l�q]��«�A����t"
���ی�s⍢x9��i+ǃ�U_(�XIK��'r������>������t�D?g�J��Q�QeWaD�Z�`r��� 
f��A�.D͐���~�v�T%���O����!��5T��j�^�Am5����[��o��w���)O�T�`�����k11��f �/Ǐ������wP�D˸I���Hpư.6@;e�ev^Ta�rpPL����?$��^��|���!I��{�I6�&�Ҍ��糠9����b��	�d�����1]�cRJ	i��T�
}_2�q3)�����x#H�^'��|R�J�[Ho%�ք_�����:B]#���R�&��w�h8�8��I��� ��Kڻ�t��^3cZ�ދ=֬n��lt�j-j�p�ܾ�Y��,I����Q�^C�o.B��q�ְ��2�s�n�8�}������4�,/]�e����3R�Qq[�{�ya�t��Vh7A�OÝ&�>rb:@' ��D9�K�i����[�>-S���v�p}�Ӵh��-Qf,��=8��d�o��(R��6<�;!�dK�����L���@d���Ʉ/k�:�(�K-;�T�m̊���p5U)-6F���������i�Y3���ؿ�me������W�8����(T��E�����������&����xRK�����Vj+��n��>���EY� L'*e�Ыj���$��R�+�J�5�a�����sH�����C�.�����h��k��Ҝ������!��"�fR�X�,{�+�*�̰0D�i�sPO�I g�+�`Z�i�y��HXq�!∋@��g3h~���;���b�M����n~;�W��M���ٓN��5*y��Vu��>\TRv@~h:7h�}��)	��ۧ��Ar6�Y�a�T�!Ꙙ�����_%G�OQ3���bd�.�-�1�"�_�^)MP�sS�|6	<���~e��B6_��ؤ�[�ؔH�p����.�x�OMQ~qA۫xF��#`@����T�BK�\�*���7�8�#��aX˩WTj��uܸ�*�д>�n��mI�d��ߎ����s�*�����T�qo��s���nܶ�Ƚ#8z�ސ��0����҂g��j��R�mE��ϑb�3���d������C������B�m�<LN�m{�TF���*O�Q?��̬[y��1���7�����9V=�[�z�tudh药,�@��X;����k�x��(�����/V�!V�����Ԕ!޾�/�k"Hd��jl{�p)�k�@mh�p{�n�p�����W�t�	3����c�zkO!"�gA,���$v����8���r���.���kf�����
lPN[X�!�������K?~�m��i.J�C���Tĳ<9պF�"�o��5��N�z$vP-v��N<��,�mL��k�Q�ĉ��Y��So����+�ٍX�������#	���*h���d
��ܥ�Kh$��y	8�d.��4��eA"��,a�&BG'/-(���KPg�!��Y�:�8��� w��s�sw΋�q�,IЁ�c߮?9���Y����~�v���#������c�������f� � 2ޕb���`>�d���-߃� �+�
���aG��1��Ɔ4@Z�U󕸒1�-x-HϨ4��Rr�3Rf"��Xi�E_��Na8j�q��|�U�7�܁O&�����v����։٦�ix��?�9V�pЭ��(`W�G�c:���^޸�#���ʍavsjj��t�A�ԱaNf�AO��+�Lw�3��pt�7�[�QԖ�6�l����ڻ>��A4�my�g�i�x����KR�1�Ŏ0[v�0sǲ��"��'�;X�t����)U<綆S%�LZ����_ׁ�<5$�;{a4؆hѳ�⎅L~�է��F���� �Ӂ<!X�3�^}�#3Z���P�b�kܻ&b�[#٫���d�Q9W�3qO�0�q��,-h�h��s�ݐ����(��-�~0H[,�Xy�6){F ��?�?��4e�6X�����1����l��hRl�õP&#S}.Pv,vK!t6�:�����utJ	��`�'�(��Hm���w���l�`�����-K�Y�Z�0D0�4���~�%}�7gO����T `5l=���1#?��V�;~J��F�kH2�^j��mt���hLv��벥n�\���@W�tռ����������n�(r|�mJz���/�<Z�J3�$��I�W����n삗�N	AX�a���*��^~�O�l�c����<�@7C��ʃyM�ʮ�fpH1r�[�^v�B��2�B5^�
���e��\J2}� �����=b�쌻���Y.zc{i��8"eò������~���|d����1KG|���{M28�l�R�b2�z"�?kRpk>:���!�N�+U�I��=�s��pNI���o�����yTu�P���֨'�F'�.����Ax	Q%l�3PI�!ǘL.[9+[����5��gYt�i�(7f��_�*�������M�@H��p+�����HQ�����BF��Rm����&��;������� y�'�#�o|�P&��2�*����<l���Qޞ�l��C�'��X��@v?�D��!%e�6�/�g��g���QO?��-�&+WM�	���,�w¢���#�o:�Zo�F~'d�4� �~�u��r���cl���Q���O�"�����M�]�e.ƭs�[��'��c���F�j�w�-Z��B�d�)��'�vF�mo%ᢎэ�z-�j�X%rf���]����>��9+Hoo.�%Gr;�R���6��e��5h�S�w��	R/ǖQ����	Ƽ�[8�A4�]w.Y�qɓ�P��pW�
���:�f�����S��:������ ��vV=�Hʇ�&��i�B���R��R'l�)&D�A�6C��Ǳ%�*{(�@��Ϸ����|�A=:A~�^�+���@�O���u=���RKL�@�5)H�l��iY3Z
�B�{� ��y�\^���-e�'ڔ6%��c�>^x����PU*_�����ϙ9�g��3��Z�{�E�җ]|�A��G�Z��=$�*Յ��i��J�����;#��f���1~����,C��������1�sE��y�ɫ��f)g��1�V���0����K��ն�k���+��7^>i��H�u��4�o_��"��I]\��Uo}��7��v&�u{cT:�j�Jyc�%hlSR��ag� �l�T:0��I{�	��1bOIp�SDJ�?2lH�7P��C����Kj�6��(�!Ț�',�j<�q���A�3DEl<6��z7;kc_�l �⻷��1�xW�R�ͳI�E:��Q��\H�rJ,���l�
)(�O=h��8���{�$��k�4ۘ_�X�1l�g�J�cG��5*8
#kN�>S�g�o�%��������U�Ұ���N�̷��\i�|�Zى��y8��U�	y���_�$�4��v�z��?��pg��Q�~��Ѥh�A����p{�h�g��cT�ڙ�M����ɬ�+�Y�H1�2�膤b���-P��VRi�祰�B{�︤�]�b���ja��%��U��~S���*��* ��)~sXb���C�o{?-C$��L*F��^�<�3��ٵ�0�0㢉n��$=NC.�����W���0!��*���]f�e�llj	��4�p�i�:f�T�eI��py�a�q�P���x��Jp�ên+Ȥ�{�G� �F�]T)&�m�Ҡ(�X��|���q�b�I��p��Y4����<N�ܲ�_(�M���n'A@�ZF-��Pg�DU^uUeC�Z��JȽ�1�����	e���y:&ݰO/X� ��$h��N�L/��d[�w_񼝱P��\_^�a�^kp�"���dc��v*�śż��E�r����g`���Ƶ���A�,� k���<y�)��4d�B�Px���Nw��aW���E�p�S�7o�wvyAi�6��>���ŷ1-�G�&	����I���0)��Ar�j�%��О�������Y�N��j��y��Z�p�@c�x�؄Ծ�~�����
�f�W݁�44
e�3����m)놳��x�9����AY78��H���^H/`>}h�r��y����o�ݲ���7R�XhE=�@
����R�V�|NE�
䅑�/~�V>n&�Ru�x@n�H�V����>�?�q���l��� �?�3��(��.A�M��P�}� ����;����.<�w�"/�o�= �f:0�3��0��w@g����Imz��1br���7���G`�FNg���m��3oe2��L�*�IG�X�I�~��v��E����9N$�K��pk�A|�©)���x�m
	�<T,�7���Ǫ�FC|�}� �AX�[�!���K|8��> ��-�8|��t$H<+=<��t��!�h���"�ZJ�� [����Ydϊ��2j����@�}L�䪾��>j�S�ս�����3 �%�=�`K� y�9����ޔ*z ��|Un)���	~B�6JZd�7�ф��-��H=���Ҫx��RmYJ���E�ؗ������<�,�듸�}.��������jS�M��|{�ۑ,�����L*��hhed�P�==���nT���u�g�r]��Ep+a�(6��)����_	�G"�=GZ����U)pj����d��I|i��O�(`d��0�٫m�qUa��K����|g�,�f�F�k�$+4��O���ڭ�]�VN �JB�s�cέ�J�@���d� � ��6�]1����̦�}J��JR%��?��iг܂��^�-1Kw�����-�����7���2p��g��aQ'Ao�:�a�ۍ�� �e�s�y�����Yܥ������|j��9B��(&»�M�"\fEfͤ��P���8��~U�ۏ�m���IX�m���&�Nf��ͭ�3L���%�:(��L���&�g��Jnی��C�v������-���r������]v4Yй�k�x��J�I��ti|#p)ID-<
<���>/#�*�M��@�v�NAv�$U����>���7�v�x,�҂9�T����7�8������*<d�ᗚ��-� ���}�L����S-�{J�9�0[��8�2�o��� �_��5�'h��kBnٕ���?;��5�B��\�ޱ޽�o*��Y��F�B�U��
�{ؤ'9i�:.�P�hB,�vi% 5�Pi���aм?a/��vA9}���dz���\���'A`�AH��F�,f^_4�Z����f�%Mk�o�Gtz]�V�v�r�v��W

We��ϭ�&W�R�b��O�n*|`Z�`l720s�o�M�A���ytÁ�*V�R�Uk��:6B�lL��3r�����@/'�Wә�U^^'��28�:�s�︔����9PԾ�U�M�d܍)�� �fcF�u��w9
t��~大�@coz:�>�L�<�� @y޸�j*�����4~��,b�]@^�㚲����_��}k[�F.�з �<���.�Kі�#��<+ <կ.ZM�35�}Q����k�V�*�Q�5��kC�d�|ٸ\�	#��]����Ғm����d��R�>f����o�8��_�1��RM�����j"���/�mR��.��7U��g#�;���T�X�<��֐zy�-@�_�ŷ�l�� y�\cm��c%�(�Z
�1С�� �"��h�ޛ<����'1�7�y��M�Ε���Ϻ���F�sA�6�\P����<S�7�ׅ�mD�̃��QpP��0 �502�+j�=w�N��Z1� �E&��dh۳�zˉ"<�R?%S	 ���!�|�
�!?kb��
:rT��r�SWp��X9��=���Z[ºt��"�K�7�K�=Q`9+� �:`8�%;S9X�<<g+rK(�, �o��������Lb��s� �\ƅ�nN<}:�˂ͫ��׊g\m��)[2�?�0��c�����7" �b̘���k-����Dz�3z��9��ꗇV�%t�h���Ӄ}'箐��L7�({`�����8@:e�`��ů@��* �I���_�����<^��x���R@u|�� �4�IڶNol�iB ����C��ݨ�.Ȇ��$*��������l��y���:l�v��C���Tt~�6ٻGT7!g��]P%�'�S�N��(�2�0bf�.�lK���Ŏ�[�A��A(��a���9n��<B�$Dw��Ԫ4,�{��t��IJK&���F!U���^~�JzRJ�0E�IDu�a�0y����D'��6��mK,��jsE`���]��&TIH#t�G����+�v���W�G:H3��*�:�B�q�D5;�#��w0R��
y�"% I܂�"<�oU.�ľރ�L��H�Bd'+}��\�7S�)>"�PS��0Q���{T|Z����ap*�Q��;n�(�3dm�𩖮v�q�|c�j{�1C��!AU�YEZ"�O��$u}�GO7��3�m`<
�oް���)���	�J^�7U��Z�D�Z��fr�-�]��UOTQ�7�ͮk��ɏ������o��U#������в'D�(W�3��z*p��PA¯�hnW���G�n@�S�U �E*��_���xp��1���9���2+W> �����^��+��J�\�b��	���o�����n�(�4�\v��ąi�j͕_�͆!|t������0�j]_tO��n�P�`�1J�ð���Ip���H;b_.s��!+fhQ���B7�-����<ZQ��B8%�l�E��z�sW,�+v_�R�DS� M�/r��e�$(��	ZUz��~�R%�hb ���E�e���پ�)~�h���ln�\rɏw$J�K�%���~t������׬��Ș$D6ӝ��@��=r��48e �v}�P�99���#
C70��1��a�1X�n�eF��'��޷��y��)kڸ«RyK�>Pd���p~�3�T�G/a�خbj 粽t�]�(`�W������y =����{�$����FX��_疤����c�u��n	�$X�����=�D���J�f9�(��F? ���
�J`��VJ��=�oڐ����w���PO������qY_F�9��D8�U�:�460��d�)�E��>(������.�.�N�f��nm�-PQ�����k��|l��$	P�b��3�5\��,� C�!���D�?���ޭ\�͔��|/�r����J�]A���In�+�n�_j�7>�Z��P�$��Gk�j'��S�>=�;� "">:V�~�AhL�H�6f�ʡd���J�eٞVǔ�(S��5+��f�#БЍJ\��űU�1��%͟����k#~N�7Gю]K�Q��b*�-2Z�ߪ��<��7���Sp�5�(��]� ���B^Zf���&r+2���v��fv���K�9/�{�2�a����j�K��Lc�}N$&Vʽ�I�?����[-�H�:s2�9�_X�-��nw/p0�ϵXp��d�m�Z@�ɻ�L��o�7�,,K�w
o�\�G�sV��=�����BV��SC�>0�[���`�Y֮
�����V�n�N��q���*�l����َ12���ݶ�I�#j��3E�����qm�<��[������nE�.�<�Y���lSC�h��-pG�X؍�n$�6Q4�p�������!��4�T�{����!�o.�˞�8�}�HfVv��y�(�� �z�8�ƥ;ȴ���|��hW�|%AP>�o09��癘g�,oc�)oL���I�r+P�
�7_=�y�Ůى�+��_�)�D�f�p�p�*A�B��9���$f%�-΋w� ��Bn�Ȟ�crI�1�ţ�����u�34�v��膿C6d�)4
9a֗�A�0?Eb� ��g�P�#Z�kR�e7��w�u꯴$Z�C�xǬxz�<O$�n�q�7�6p���v������P��qf"�nľ����V'Y֊����Y|�Zf�V��=ߌۈ��W���1���A\�qezc��l����$�*�e/�^aA[X��huв*��=mH�Ġ
Djw�W��5���Qrd���1���ܱ^(�g�c�^rE/ŭ�h�	�hf�s�`+�3��.	�8�Z*�|PҦ�.1V��p�[xȿ�<�8&.iaf�[�3��9�,pf!������^ؘ"�T���������l0�*���/u�����O�t���!A����Y�I�9��6��ޱ]�_&{'V&l�۪h������y���I�-�3!�vIU�����1ΰ[�p}Ů���9�9�den�*.�$s-H!�5����?�ؑ��
�������>�(��M�y����0P�.�!\��{�[)3�]�q�ݾI�sa̧w�bKgK���8P�m�P���.$M⦔��c ]�k��f��軪+�l��T����Q�?�)���Sk���7D���׵����3V^�d�Լ���SÐu)21m��ǝ�L�I�ޡ ��%��h?��W��el�H�<6��9]ye�S�Q����j�4��M#�X@"s)?�؃��0�iB��ɠ�onq�� ا��=�������{���2��ί'[��3z�@�{�-8�c�0�Լ�J��U��5�r]�{!�Jɨ�0��#D�q��#��"�0��mV��'q|��ȇE�b��c�W�����j��̬E�wa�bP�yd�Wa\��x�?�*��2ۅ�h&�����<��3����ܽ��H�׈��%.`��%Rg��gnI<��qx
j��=� ^n�����y�_H&e$l��~�O�`���&GM� &�e�5&,g�*�g���1�G��d�R���YϦw;"��w)��hX��i�M���<�<o*�@a֟��D�(hx�"\�J*�½B�P,y�Va�t�N�S�~��27�!��[1 ���˺�`T����E�Z��b]��ۂxk��K� uQƍ������
̬
��rn1֜
�mukpG"[w�P�a.�FߛL�yLRb�h�!h�hݥ�J����!�<)��f�;	��h�|1��{|�#�b����8�[|������j���7�?�������B�|�8l2�W�_�	��G������G�Ѥ���3Eڐ��<�xw6J�w�h%��%{��TE���oAk>ϡQ�������28��9s�D�i�(7	%n0	��˵�g~���҅l� �g��$v)Q�qV�{ͧ:	Q�����"�pL��P9�//���6!8L���z����;��P0W��x��cm[\'�0�����02m�臼'��B�n�ce�s��2"XtdAj؞�KS�}��Z���d�����R���a_1��,�'l%�)Z�Y"��,x"D���}��OI%�c��|��s/��7%y�[̝��1~+�/^ߞf�G��׏����٭W���BQ[*���~ᱴ�6H
�(ԞD��[���࿸ڐk�z@�j�_���@ �����-��_,/�rS����SE���_*Uv�R<1	!lRS�O�=zP���_8?|s]�����?����z��/���f�/h��&$�F`��hE�x�t�*J ��`�zX<g�0�R��7��}!b��tp�E�f4��$@��3"Vh��ޟ��&>yMY(i����IV)��3.�]�G6q��OV��x=�� �2�?+\�5�Wg�_���Ǚ=. ��"�n X�ŭx�L02�
O�f}��c�b�L����q'�0#�cc�?I�4������4�`۹4~ M��ZW�C� y���}Wms�\���-=p��:@'�##��C
�"X����e;XG4�HϮ�ctΉ�5��͏y�>����{�`M��ktU���}��pw~de���H=�%}��?[��u������]	`o��/� ��M��ǯx*3���Y=��\�l�v����X���M�l�������j��kK.�e@�z��RP��Df ��'DO,q�(�8��DKK�W��Ke� u^�_�p���P�Ɗ��%I���P���]��8��eG��"��o	'eg������u�����o@�&}��g��t�TG`I���T���\�ޑ�xAY���I���"�Dw�-�1� rњg�6�5�5k�v�0
%�u!�[�Sl�"��g��%�'מ�.��^2�
/t���nC�/pu��	bq��`�\T�A�Bh�� ���_!��Z�t���3�֞�)ā�~�l��}��P�0��"�X�"���o��'�1��,������`����-�k�qL�YQ��mr2�y�1`�pc�,cb�D�ϔ�+Cu�[2I��/�����4���0�Q�i-y3�ܠP �V�Ndw�i_[kq%��o{���Vk�l�fy�ct�$����ob��	Pb�%"������dQ��苨�轛��B��5���bk8����d[�*��%(�5��!6.��Ɯ���B�C�̃���4��jŌǲ��Ց+����N����^�j�Yт+�n�x���h�3�-�p��>wz��@aX�VrU������A�&�s�ujm��Ƨ���#h,30ֲH�V�|n�ꥍ2]�L��,\*�3+���r6��'�dBA�{�I��0RF
���UoG�bE������T��r�<0�S���N����(���ȑ��ֽ�A1l�U��	w��ϝV��d�y�%==�옔#�Q�������%���\Ki5�
�9�wZ	��+�vN�?r��=,����1�v�3�y��5YK��(��+��Y����(�p$�dF�Z�+T]�{�Dy�	vO�p�x8
�~HG��6�H3Z�����y�?'�9K�;�%��T��jo8��'���UX��o�A|"�i�mO2��u��Q?
9۩T�˶*)�g���@?��塗������n�\}.���.�q����;:K��L�&vG��]l�U� p����aG��Q��y	v`I"�[��O���wς �`�aLcb4��ԣak:9�?l��h]t��~=2B�ײ$|k\�D*r���/�I"�Y�%���	��\�C�ٞ�(*.�Mh;��yC;5�S�٩��2��6^eY��^�(E`��6��z ��dz��?�^(5
f����$�A8~'ʨG�mҵ�͒O\#�e2��e�A�4�3�e����#���g���c��-/t�#q������/�O
a�����9���hS	])�19�C[���$���G-oQ��Ju�*��y�����$�@���ߚ��������'�1�+XԆ=���)����$�fHp�@x�1�aݮޥ�]ޭG@�[�7i 廋K���͜�(΋lo�2���%�&��Ϯ>��7���G�ăb:�#yTʇ��
��I������Gі=o�T:�]����HPf"�O=�Ǿ�3Po�[��<�k�����~5]C�������J��X2Lڀ9�H%`6�N�pV~vQ0���$�؂���+����E��A��C�l^c���f+��7FJ�	�>� ��)nں��KȻ|4s���8��A�`��u����B6,�.�V�do9��\J'Pԯu�[�諄2�n��N�m�������qH��
<z�5	�gk�¢�����f2׵����=��K��н�kSN��=���
�~Z"6d�# �ђ�ͱԂz���f�#�i���qC�z"�a�s�}Y���BƜ:x6J��B|�Om,	���}\��z�t$�䂶S�z�UJ�߰\�-����&%V��as�X�(�D!�<9�^�a�}����t�����>!�4/��n�Y!��-1]��SUk�/�r}��o��#q9\C�M�zQ>;M�h2����>y��������ŕH�<���g8���F	[i��1��ȥ����x���6�Ȋ֮"xs(m,���m�8�����]4M9�٥ Љ�Ƈ.�	��%fR4]��*��eu���n��aQ�v�O�7~2�����^~�奷���]`�C��5(C���\��_C��W���]\{���Hװ�uf�}�I¡����
V�����}ѕHh����w:d�bzhLhSE@��:W����B�1����/�'|׌�6@t�������	�ߴ��!luт��oκ���V�h�0Vժ�*��72��I*4���$^fh)8��T���:	�p��Uon�a��R��;W�?�K= DA�D�6	�T�.�����1ֆ�@@�_��s`x=��R��%�ޒ�0���q���ѕ�}�F�6G"�A��u`L�M�;΂|�P�P{�9W��)��;��Ŝ�^��<w�{�VSz���)��J�F�#B���,�4�=��m}�'�e2%O�YGPf-�0�8&4_�R�>�ys���
�ݑL�	=���Ag�\�2?���?}�K�Ac95H3�2}����7y��9���g��&B_{�`O�	��\r7.+��H^�4\�Es��������Z����Ĕr��J��e�&5��p���Q�k/m�J@|{��f���v�^Cҙ�9[��8e<�$�?�M���!ܑ�[r�fœ_mHa����"$[����p|�^�G�	�`��#{��g3NL��FB/���QF��B/"��2�8O������� �稫8�:A�m���_��z5��\'�LA�8]F� h[DČ��`���R�ꨨ���Jk��G1�-��K8�R.�ܵ`!�o{6�k�;D�� &�ҽF�v�TօpZ?��>��$�7�����=�)�u���ǆ�e}�J�Gf���X��	T�%���.C+��q��"�΍ �8����l7�:7�LQeM�9�H���{\��)51L�IP�O��������d���h���%,7A��Ɂm��W�` �x_ Z��$��@U�����ԤKVjsB��m��$�2R���E^Ŵ3�!�p�R�;��v�rl(>\FMHH�~1�Ϫ��c�mn5�۴5PBIYCkܰ�&�2���������ƅR�����%����^C+|O�֯Nq�vO�ʏ�@#\��9���)Nj?L(��6���/nC�m�.S�:A\�rz�5l�7m��(����67����`�7U���V����ӑ�yM�|��	��1�5��'d����bav�bIBޯ@ű�x}K�E�Qe|���Y1��!�pOz5�����nņ��;0�ӧ̯�:쮮�;8�}'ُ{'��LωT�dy�������k��燡p����Z��Or�	��8�fy&��4}6KQ�o0�K5I�YB~7�01�#EM�W�an+��k���,��0� �=:$�3�ZD��AO�;l�8{��7��Y(�V�e��b"���Y�W`yh�4ɂ�|_�X�?,A� P�8�����i�Hc��̯&��BC��f�-T�>���gOju�a%>���@L�Y'k�[\r�L�Wx�;4/�u�R�ʈN��ݑ�OٜI�Ĺ@��D�����C��[�/pNǅ�og���£t����ι�_�tTt��
KzJa�t5"��������E��>��eP��p�;q�l��ܹ��]��HH{��Rz�2�D��ЁxV܏+/E�6�ڒ�7ew< �����D�����4������u���;��vk͓��ܯ�0�P�D��\�0���ݕ�)c�aH!"����P�%q�%�IH��&���me�(��)�st��(���]�����j����w��n1��uXi (*���t��-�;����N��~�#��7������?Q9EO�kRC�Rz��MK��/��,L	�Fd�+��K�ᱮ���rc��C���+���t�#���u�ųo�iÜ3�{m���X����|�Ct��
MDk�.�5L��)��'BP1���s�x,$�wD�l��8��\y���-�*X�nт��x���~]nr)q-9�(���~�w�`kn�K�&<���D0kg�a d'��ol���Dyg�^�g���ѷZ5��u&�gm���8��Ru`·a���Ԝ��& �;�`M�ߏ�id�B�`a8��x�v|��X��ر��ÀΟS���&�e�}Zƕ��B��Y$�L'n���)"{/٠�Q�t�ͧ0�����E��+޲h6L����p�N����8�8���FK/==�`s�����@���r9����*fzn�ןר셤}��q&Q�\b�mW�n�X�����W�r�Y<�f����7t`�7X�J�.�dy
@������hG���R��ҡ�9-�פ j��	��g1~W�0q'm�0�M��",{��5����ϩ̥�dD,�h�1��?6�+Wo�>�n�D{�bSU�C�O��Pܞ����P�O�ѧf
9p�y�hq�>=�/,�:V�s?�M���YG�V�6Zb�g�:jgR��^Lv <��׽*�~|���(�qE�p�r���1��VWu�^�]���6�Yb�m$[�sc��p�[F��{tp3S۾C R����"���:`b\5��۬���$��}`����˽� �����f�h�Xdſm�o��8�v�m"��Q�ܭf�F�.e��Mu�3\7���s�>e/���k�!`�U�1�E�J(��1ζ�pp���3�1�%:/���@�zQH��E.i�������8��y��U��$�*�H�~[̢��a��;:`�,qQ�LY��8�kg���S�SCg��Cu��<Q tl:��$���/p�S�ۡ��h�ŕ`��G2[��4:x��:��
��e2��K�N����.�;2�R�K�^��k*!�_瞐������6[6�˯���7f7<��_DI^CYa��/(4i���H-�*8��|�[�!Wpi߮�$7�1`%f#J����S`�ڭ��Np^�oeP7�8韮�����w��PG��;֠��M�=0W|��c�?1���o+��Mmr�ر>�I�Һ��o���=���B�B�RfP"pOqE��-�=����v��$��K�*�yH#������&�TVIƎ8�м�c�%L?�m��MAk����u��_���)��������S�e?�[ϐ���80z���*���g e����G���?	�˹�F��Y�
�Ǵ: �eL�9�����~��l:~т�_X0�u�m`m�W����h&�@�!*@YZ�7���8dL���B�[�B��.C����;.��w7�� ��{ԃ��#�n���/�竝�����%Uՠ��:��b����]韋�����=6��J�Ч�{�T���X�9�痠p���W	7K���܆�.��!�wd�vn@�Ȼ�7�Fj��Xn.�Ws'�h�f����D��i�E7QrI��)	}g��jh� ��yDXYG�7�°>��r���/�Qv���gw���.�,:1:�����U/��Ic���i����O�~|�?5z��~?B%�e���~��^'eq��jjl�`�Ն����!�f'����A���2aX�F7ʴ%���S$�Y�}�v<H#|P���*�2Ұl����>j�J�Ւ�L1�(�x$���^��y���A�����$�=����SILd�����N�3] �P,�AA@*���D;�r�^�8���&��BӋi���U���W@�44�E"�$(@�f�i�.�0�8:�7��_Ӽ7V/�S���*�L#�؎eM��é�k~�S/=P>Kn�0��.cy��Y\�c��I��=R�e&8kky�J�|kȯ��Y�t�}gP��v���N��@a�I�7�B�Eڟq����	Q��&��`�0L� 	}J���  �!��P��	6#�/j�	тC����H��{�;s:E8b~3��Г���V �H���/'�O�G-�0	f:F\1�\Һ.T��t�غJ���ހ���R�O,o}����z��X�S�}�����/�<��/m2��yI*ٹ%29pR�.�����5����f�;`h34BF����C��!M(�!aw �[@1bŮƖ�aĴ2kD��8�%l�'�������_\M�'QJ6ަYi�$"lG�
���'�m˥+45��.�&��p�!ݿӰ;"eޠ;--���5`D^��W���J���S�g�&��o�̢�t�����&������"<�g�����r�P�v$)-֜@�L�@4L�������.��68�ʿ6>�8
y���Df-���qp����/.X��]�J���nC����}�f�`�"ް����c	oW�=#[��R�WǾ���~`��-���n7��qy����:��]k�U��4^�cz�g �bZja�{���}���W%��#�p���%kb+�B�R��2�xG��y�z��e��|�^pL�%�ҀjQ��ֱ_��Z{�4�;�PeG|�����ǯ�� Aͩm*1�Y?��blSߟ�N�ΥQ��ڧ�M��8�M����P/�P8��z�˦`�H9e	sӄ}��;{���^���7�S��n/�a)R X��OxT�v��;-�}'f�`D�";	�	��Gnw�#QRt}9;h�3w�6��֛����?L3�:k���5���#�e{�/�٬sh\����sr��_��k���%��ճ/�bMMƩ���UI�$���J���p���K�p���CϨ4�����mBp�i��iD<� �r7n�K/�m��1�|�k8������p�M��l�X��j�,�ʅ�?I�lrqr2�^����$�3��?���Pήv0>oS\���F15f�n��A�h�G�>L�-,��j��������K�N�f��v�w�ҭ�$>��sv_��<D�]�����.����\mJ����$��������&��H��t0����N���m��aK�#!�i��j�m|=a����U�tӚ;{ b�Hj�i��|���ݚ؟��ise��R���A�/� �a��j_�`M;�Rf3�pb��J�K�g���������AJ�����Ӈ8C�Rꚷ���[����X����+�������� '���UXs%��"P(и���ʪ�bG�$�q� \��n�`����(#���=���@9�*��D.��Ѳ�OdEےH1r�^�	���Q%���+봌��%%W�'+�m��������&��^Q�*�j��qk��]�Wa�ZT���1|2K�:��O5�1 >��}Y��O�,�`� �*^/P��j��X��8��n�'��t��G,<9���~e�7�h�;�u m6�������%MFHPef,�Yl��(&�QU}��B�0�X.R���3,�B�fBk��H9O gυ8/���J��l�\br�������'&���i�Z��M����!�s��*�}F��&�5r'#>�,PL�Z��f\c."�TK�jwӛ��.ME]�[z��� �[�Su��f8EB`��*�������M�J�3�To��2�c�����<�b>�@����h��vaګ.�/%+5�DH8�k;���d�al��]�6�Okn-�/�����5�b�E/���O��;?֭�A������1${���$/w��ܪ\��	m6��m)*���JL�b�Ht�|4�,�M�nL���`�{�{as�S�8z'��E�U�mD�2�:p��|'j@�Þ'I1����:���=���� ��f1l�s8�]+q57�Uk�M��@�/�M�j/ƃ�6ޒ��J�lճF��괛��p�a)�'ۡ�Y�X� �� Vp�����扤5{,�v�T�+�8q�̼h�lڗTr�(kY��MWe.N ��f�w/�P�B5v��n��F�j��i�r�p�G�P��v.K1��|ݱ���[����P�k��ݟ`��s�g� n̐0�o/B`�Ub2Z]�߿���^����.���@�;���J�V5W�*�}H�K��}�y��^%%POaF�t���T���sc�#�0~�B��p$� �$�g �rpL"t��Ɉ�w�������z,��P0VW.�ܨr�]�|U�'�Ö�'��)����s��We2 O���Ey�x�C-��Ә���fR�%�ps�.�<Md��w��-�%������h���;��!�.e�#0�)ぁ2�h���6�K/���@=��ݢ{��VM����7Y-@45N�����#�iuB�Q�2�d�"�M��LF���A�x��k�M�7���+�_��:�V�e� ��i'v`|9�Ikv�Vrqq$���T��1�=�iT���&�:�t�Ĩ"��7���?zNVi���m�����}��pZ��\���ڹ��3����K�}��x��1�$0Et_c�Yȸ�`
r��1:x���߫���M�ӎGޡ�������{�1Y4}���D��2ץ�a,(�}DC�W�������<k�SYԨ�5u����c�0�??�������-~o(r���Y�My�Y]�����̌�&�( �����c�7�a\B�W�z��!�<M����hE#���6F��P�^�>�S�`7.Σ9:uYL	�4��,:-��&�ܚ��ƽ�!8gp����>�ő*�z�f#3�YN֮�����m����s�q]��fւ1�`ŹEܙ:��d��X��mΕ2�OHIX���F��5X�f�"�{9mY�Q6�ᥴ���J�ņ����tb�ͶO��.���ru�:)�a�oi�%���ע�N���JН�
�m�e���C*HX� ��y'7:X�>�i��g�1���>ݲw��9klP����yKnΫwq6�ת��RC����|�cQ�C�X��!����Mk(���-���s�@1�J�\ޚ�W��B�{�ˠG:Le˰wB�C���&l�_Ub���t>8����Z��4�{&,
��;�N6if|��5{JLl���wԝ���J���V��G���� ��:��	5���H��U����֡*.�v��	;��Rv��D������l}�H:iT�cW�'���S��dJ�s��O3��[᝽�ү3�jI{Z޳��~�c��ɿi8�p��"��bJQ����%�u��
a����|�KS�Ei���{0��F�ʖ]XUZ��%Z�� �6�I�1�fd��pY�\��G�G���yk�%
ܠ�qx�}^�^JX�k���b6�Z�壤Z�z.��ʐT&E}ҽ=Ee��M9�N�3IG9��Ԉ��s���
-G7���!-P��p�������3��+�#r�}����_�n�I��p��4�S�0jLR�D�}��s�F�WE�G�jC�o���N՘�Q�� ��N9���U��k��l�D$�l$}�ry7X�Iy/td�Q�]p�*�	������ �b�V��|y^��Pf��L���f���k���m�mS�4I6�,&���������=�O~0�b�z�>F4gf@1�wza8�FXT �����hCvs��yA�'E��c�0>�	)3N�8�b.�.Z��^����F��k;_4z��e`���t3��1�����&��/�^$�*���W:�;P���IQ�z�[���,Em�R�0�~�����Jt������	�:�����[���i~��T"��ݏ}.F��x�i>y	��ð8X
�Bfh� �T��8Y��i��B'��]B��ju�}�'�������<E��fU=t"��4~Iq��Yn�������d:������U/�w��c[�ӳ�l/�)����`�?���6�:=֬&�fY�Rз/b�3c�71d�R�rT�H�Y� rZ�@ϑ�D�6e�#C�%>§��0u�|�	��[WE,�#��|D���<�!w�̠!Ľ�gM+�R�5��9�g��c3�[u"�Q­1ݩp.�>��y��n���rai�Ln�7�b��;�J 󜁼r�-�.G���V���F(�����3#THuzs$].o,JǍҘ���_��II�u����Q�Y�7:40�Z����V�`w`�F�}�����\�M�J�]_	��5��aC0[{*dDhB���������* �r,O�>�-�1p+��u��뷾L=|P3����ds�p�G{��a1ת~�v�#��*al��<YHF�@���֛�n����T���4�M����b�H�x!��1G���e��`�&|�^�b9p�A��[���4�2��:>�H���A���ug�ɻ�矩MMUW�`��R����H�>=�Щ��S����{�"e����]#L!�n=�)y^���\�*�Ɛ!�u�M"`=��9�]cH؎��o(J�B�����^��Nl
�Jn����1�H~l�E s����㼭j�.���?��3 �WZ?�H������Z_6��l�B�F�(�t-_d�U6lzZ�{�a<��0S�W1��&:�J��fg���o¢���b�/Ȕxұ�	$:t����ă��Y*%�Yڌ(�w��c拢XT�Å�󽅗z�N�}�Q4�w�]�r�AF�B8XE��hęxؕ��o�L��f(#��8�?H�+����Z�(5
�݂e6^��e��L����|4�\�_c��/�r�xi����!��>�k��p�"�2����fk^������C\:�
���n�S�b*��&��Ұפ��H�pgL*�'�YbJ�4ήf�@Ƌ��M���:Ϯ��s|�y�}�T=r]���Z��㤛a:>�-I��Ȓ�ؘY�I}�U�>��W���R��"I�Z~��`T�L��[6|Iň7F�Xmo�Q�����to�k�����'Xy���u"�W=ZzH�>l�߰�6�?E�����!TW[j���ɸ�l����4���c�\��k��ü��V3�qֻ��gd��'�9�PU6ӡ��zLH�C�Z�F�Vx�,�D��;�W�y�H5z��R�±6��/���u�
�d��Kv��7�6�,#5[w:T�������i�H�[^�Z&b��]�}�0Pr�i����II#_�y�+�q		��߼��� �W	H[u7���į��&��XFL�*��n�d\�}:%�H���]X�q�z!�v,��m���}�1bk�S�9��~�ǯeI��C�{��]B���Ȣ`�)�[�伥�R��u�����O*������w8�~���PD�޼H��n�:Ij�Ũ�p(�i���O�}�k΁�v!s���?��׫оX���V0�o>���P9v{���9m��ԅ�Yp�J��A���Nu�"|!��Oo	>4f�K�ɛ� ��p'h#Ս3Z^:��t>��;ʮ���<�������|o�$:�����! ��君 �/PXm�e��-���܊%��5�=C�-F�ŕ�zq����9����m/�@j��NE���̢Zu�/� !V�U�E�d��M���?a��������i;�!��Į����j��*<� ��P��_�ɨ�g;��cͪ��e����H�vIő�3K-s|5�ul��Y�~k�Dk/�2���� ]%�Nji��;j��B�R���:1~˕�=U�B-��r(���n%d�)R����XV+r�58�6߰�v�e�c���a��}3-�%g��o��_�D	 �x8�Ꮬ�6#΂쵰y���sA�}��1���h���f���\G(��k��3؝Z�&�GJ:=H��m��Ο7Y�rV��T����0?�����ɜ,Y�`��!�S�D���m͕��)��
����f�K���	ޣ�	�y{Ö,]zfb�{ȿ7ꡃr�4L'�f6�I.{�'}��+6�^Ij��f� �;���r8��d�Yș%�H���ue!���0Gw�{'_��x�������� 3�*89���BF{x����@q���F̤P�N�:��I(�%_�p�<L�T�Lt3����9�C�Ť�}>ͼǵ8�׬l�}B	nJ������V|��p�����n�|ߏ�,��-��9a�"�j���1iũ�)/�<VZ�(����d�r����ya�|P��P>�CGO�b�_z1��r��M���;gw�Ym��d�z��Y�ɰjU���xv{hU5c�0�)p	g5�.��q��(��7��Z�%��7f�)�w�d�jj
�AŚ��~TD�fx-~bT�̧�v]*N���ܕ�v����JN���*��˴����4���a�m*F�A�����)�sꗋn�:t��޻�+��8�D����&z��/�D44w2��b�Ӳ��X�M��ܤ����	��[�顨ك���[���t��)�����;3��j|�ȈK�#:%y,�( :� woV��c� 1�vD4�NN�^��Z��iY������#�Ù�RϜ�EY��M~���P�A�L�:�;�68���,�K{'�v�����Y�R'|�6q�I���6�}k��k�e���@�G��3�L5Y2��]�^9*g�������tb�L�խ����ߌ@@o��U��(oP;{p.��"F�^�DnQYn7��:e�[��ߥ�W�$���񲮘�s�L�˾�	}�jtR@��Z����X[����b��2!�pM��?���?]�����`Ka�����	GTp��[
|��̚���'���z�S/z��'���^-�}�[���Tg��0	.4���a'ͦk�.�2�C
��L���w�;�*"f6��Smj������{&�*A,�c<B6��,pʊ	��Ƈ���Q�N_��̾}�e�8�i<qW��l:�_�0UP^|����]��CAZj~���\	�<�P��`a$F����$��9��!؆��=ސK���紴�p���Mq;�8��Z�.8����I��=?;�S,cCa�/�&�Vu��]UBS��mr�{�L�!vQ��nP�t��%�l�.%#�[��}iM,����~��<��ɳ
�s(�q�ȱ�<v�TO!+��!�&�hi��]%�+;�9�5j��Y�0&Yܓ���q}>Y��u�����L����^�,d���,��n�#^s�쇲��x��
�)K�-S]�@���kA��B0���E��̑���7P�I��U�*�d��=e�P/z$�ح�(R��%y�s��+[�#�=�j�������0��a+�>5U$�G������M�%�Yy�\ΝO�~ş��QD]���Bg�Cb	�@�5��R�<�(&
˧P]�׳{�Ut��yK��7ďKۡ�����hqD��w^Rj���{�tt}�IGR%��d����*d����3E��<�9��X����O�`q�u�4{Ae�KF��P��֓�]\���!���,!'e3	��g01:�w�/X�ϰ��8��v[�~!��q�S���eO��ӳ�����:0�jE�{�%�B|	�VD�vo~�LAK���^��i72+)�v�8{z9��撁�ă1�t-P3�]y��s�|�*�F��d��s��_ʞ� � -giE:g��Xf��)ц����4q�:�o5�t�^#����ȳ��4](YĻ��m1qBCVg `fLҢ��RK�iog0�J�\�Lmp��� ]W��ì��-"��1p��g\����[L��~�J�����5�yxغZq�/����N�%v
�����0�gp]"�m���x܂�x���lK� E���ы\<S�U�.0������Z^��[���:�QI�rU�R۱t*�6O���H�����;%����ʡ��\�G+6,�9�C��)Z�@�d�QBx���[������ߑ����W'��0d�����
�V���*�Z�Դ��>�X��n��$-���O\�ТU�lI�h�J��/�Ƭ��Ei��~��ڂ`������a��[YT��vϵ��x��K��w�\�j�E�B�O@�y��zy*��D��%�l���Mm@LWpL�m��c� ��^[Tن��Z]xk,PM���)j��Y�$sl�#� m��q��G,Ql֤31ݙ�sxw;
�E����!h�Ov���;ϐ��@P�5�{m����{��]>��~ԧ��5/cD�
�yZ�P�hX���o�dz������KZE<��m�vCGv�]=�p4N^����$(�I�sVc����nJ뎰S�-+x�q��3�`��O�K�A��G����{��w�C��<odr�Uk5���^0:�ږ�h'.�;�fcDnuO�@ΰ���3�'/�M�$��j6-82�s�(�=o7l��}YT��E�]�2�������QA���7ۢ��X��T�H��v�8������_�(��E�I���N.��#�}g�� ��2�@�<*��u�����ăW���̪��Ɱb	Ris�c��L*%T��ƎɌ�§��4�����,��4�TϨh��/T��a��i�qq�ջ���D
�'K���������̔`�������@o|�����j�P�~�8�M�u^��2�h�k�WpZ4�m�nX�����s�1p&�Β�/2�]���:BND,��IAlQ^��?@ط�v4�vhV�.���zآ�{��Tb�y�@�xqY�寐��@�A���;.�p!�v�-�:�>�����~H��R�����O~�i��}�+-�w7�����%�L�3���oв�[��e(%5��Q���,�m�F����R`�YQF\e���u��-I�8�m����b<�ɥN
F{r�n�~���Wᾖ�IյQd��� �Y�)�����b�k�y��E�{�u�����m��6 3Z��󭨱n<ਖ>���0��� 1N�A���S��U$����"+���Y���7���2���Y�u��x����M�\�W^s8�0u��,�E/Fn������A,���x�x��;Zń�故�����7�����_�⣉zɐ�}:"��~H�T��&[r��Av'k]q�]][�/�HPg$�'6a\���p��_*{�lX�BD�X�G9~=j��p�Ohw���SN
�T)6tT��G�-Ѵ͓�9���Xۡ���h�*0Ru�|M6H����~W�V��c�	��I*�u�)�B��8�0���Ia'`�'v�B-U�wC�X͇��%���V��E�vF��&��V�Zb� L�Z�E̓V���e3V�5�J�i
֣k��&����h�*TUȌG�������/F��� �^7���H_Pg�=#-5"&��u��mR��^��avY"��Xƽ���k�bh"�4C�젬�	�BvM�C�`���t�?N���ј�H��1�-���)35��gQ`���
���X�_��Y"3�A�>�ɴ�u�^p�����M;wb1
X�� ;�S�G�\�iY�HQN��nEsYwfP�D�ZC��h0E
)��"L|v6�}��-M�D��~|\E�V� �m�?�U'(�C�EJB��#��]�DEP	�qۑw�`B�o&~�՝�x���M.��2��o�U�<���.IW�ǯ�r��F��|fX��/�d{�Ս�w���҈��MM���T��>*iA���GjGKiX�m�kq���/qD����vb>!�3G%�����,��ByZ�⿊�UC�nz�9S�h>.HL�P$	B����>��B���	�Ғ�u������5�C��`�]�c��oU���I���_�*�OD*�&���'���|� 3`�͙B��� B.�K��&��>�թR�����e��,��%�yh{��6����H�P�����Me&GAF��N�@R��E�	mmYO�)�k��m��AX�*�����I�a�~�'���@���!�QI5��z�;����v"�бi�+��Z�����_V{�Ւ�:�lJ�H�z+[�o�%ܙ����Ua2Λ�9:1����N�]��{���t�(@o+��;�&1�	8\_�Oõ�q�^�1�Q������
���"�����L���J����������H+�R!����R8rq��_�Y����F�]"4��a�d�������:�j��?f���,�7���1y�&�2	�����wb4K`��ٓ,8Bڠ]�OA��Կ�� �,��Ac�7==8������x�|bq��0�K�F6��v���q��|��朕��o�ru���SK7?4�m?�.��Kd�ֻ�1wd_~Bn$�x&�;<�I��7�sP����1&��'}eKu�2*��g��i�*�#����ҕ�iˁ��?6sA�a�p�E�ry�����|zo$(܈���ǋ�m �\N(���?f$��ϡ�A���.�"�BN�{t��I	����$-��|� e4R-��B�E7��jY�=҇�<-��!�OzfM�ˌx��� dǓt5�q��a̙�Xt�2�䖵�Q͆�ffƈ��1�cϗ��it���d4�=�B4`Q�zm��"�E(t��#vM��#S[��]��S�j���*�4&�8�˸�ؿ]��<
j��(ps���D�$]?(m�].����ܾ�.�1��B�~�:�a۶huл��/8,���JʣmȂ)A��V��T���T筹ʀ�D��,3�4�$J�#P��o��ֺ�����OF����`�/����H�ںL/-F���F���0�U�Z�O�B{z��;�m"���Gmz:ä����Z��lXm�(��ה��O:Xg��zr�R"��1�2y����ZwB �[���V�ƚ#nl%l U��[�ֆQR_9=��gW!,���=]�.���ύZ����r����;ɣ+@=*M��F�����5��3�ԶU�$�ְV"�� B�7�*>G,��w4t�
�o��<Y�Ǥ��OC��2��h��'4	�4�7����ywr�#���2i�##��TW��ώ֫5ko؋��GU��8RX��&�H���?�Ex/�����E^{D��?�,�L�T�*"T�,bA�Q_�~�pna�Q�Mg�&1� �)u�6rm������ܦ��꺔�y��}�l|���Ick��������b�������=�ˠ�t���b�<x�&��`�6����R���q
�x����PU����������p����xGs��õ����`�S���`�!S� �2�7pgW���F�:X���>xc̛��.��)���`g֡079�1�j�������"�*f��#�bjY�����0D�_�R�ڤ;>�d
��U�5!ݷւ;�>�JD ~`�\�K4���/n,�޿3�G��v����l��M�V��Y}
v���	�[<N�M\�߾���A��U�'�)-����v��E���Nī�$}���ǅ��U_�:��6�k���̛=T1�D�M��I�I�/�t�����w>��4��J�FR��{�
N�a
XuRی�7೉v�7��DҲkY�iX�}�~d�G��;@z�Br"{��+9	"���_7�X�&�����$Tz�Jx���Z\���`I2e�A�ZpB�N��WV?�J��j��Њ��t�l*�Ʊ�m�FA��և��M���,d[�W�gC��V�q������}z&�@��(}���Ӎ\�db��y
.���!9�I�=-�w�x(�Gj6F^����`5iᢴ�m����ݥ����t�7�TDBk�F� Z�3:��W��c���
�z@$D�a��?;���.۔z����f�^��P�&��0��(�eU�����A$������
PR��	�|�݌����̙��pG�ʗ\B2u1笛�E�rQu^����i\�f�l���N��_�΄x�ˬ���rK��[������0Ҫ�
���)m/�=KRV�<k��$�K�ַ�gem_:1V�N6� Ѧ���E������@4z�K5k9�5���2�kB|:H̉�|��j�(��^ݷ#~������Z�0bz
P�md�$�iWݎ��>_-
πKyI���{����GZ�	)���ў�)��&������q�5�P�����<SG	RjD�;�Fv����M(��~�c���d>������\r)v�ݏ��2�,�f���?��.���{C���t����>4Ζ�D8`��a�����Q�a�bc�d4����i���5&�؛�i�mH:�B�Y�ξ�c���;2�����=V�wLy��c���w�3zT��J��B3��l�PzMsK�)����a���#F�+�&Ȇ���_"����uN,l�e��ꇷ7�����Oة���L^��r툤7GW�݉$ޗ�|�k�3��c$��j�%�-�$�% �gY�f�Y��D0v�����g:��~+��-js����_��k^�?����6�m��j�{����
U���o�5�F>�8ך!������mt�HCL�O9d3}K)�<�0Y $�t�骧�����M�u�>�t&P&���O����)�sw���mx�s7A�>�ک��6����D�Ȃ�o6DJO�]F�y
{���*L�6��\���d���q�ǫ��K�W���g�/�|��ʀ�p�)V��ڵ�đ��-�I~��� n͝�b��O�}�k2{eXExe V��2F��ݭ�3���T �֝8lg���5(Ƥ�t<]���e��u�oQ���/�TĆIbB�h�*���~�5pF����	�k��(2��!�^�Y}D�|Lc���9y��� \��>��s�s����!��iV���	%9 �(��-�(�2$�UO@aˈN-2�]���r6�kRz��'Sf�몿GT:���� �1ŷ����5�q��7�]-X?	�yD��T�"��a�_�k�ڬ�zhŊ����$��e�B�Ǖن�7�]��3�1��g�%$��1�/XD-NH�j��mhL��7"�W��^W�\͔�l�l�^%4�|͢��F[e�ߴ$���|��w��V)��:�儶$*`�5e�����;��9w�`�j[��T�]4*�G���\�S��,���(��+�K�l!"K:T���J�k��2,����l�̖�=�-5I~ġ��bB���4e�{ �~�b�ŧ�raQ,�$&��l��7u���B����RԜ��2��C?�����ߌ�E3�;�-5�B� &�~B@��T �@k%���E{7��}�C	8���e�nM59�N���oJF�0,��Zo4!���!	�m�-&�Ë�fO����2S=ӿ��J��3m1�)��!*2"t�H������#����t�ӳ��_,�����4`ي�oqka�ό����3)r<e��X��8�IV��$/�v�(>�?R�ʤ�x��#�G���:L4�S"]<�V����H�+��ɢ�Sf�����N7�ИF[�����\7��^����7�w��MŒ�j^���	[���C,��
��%��߹+�I�%٦�[.QG!��,��ml��>S�v:��wj��b��$>w!r��ƴT`x�V~�v�1�@܁��<H�����y�0XFP��m!�3kjB)�U��ͣ��A���w��P�^��;H�{���r2��=����{�%_W`-��t>�H&a��������;��Uq:�3g�%����O��E�����v#2�5�*=�R^�Њ����?�mU��6���33*~}��H�}ſV4��rVrrw���&����oY��� ��^5��D;�l�bu�&�uP�F��/UU%���
?U�ˡ�q�󜍛9��ϕ1U$5nTk����7���`ۇqxQ&8�E"�p6�Y����N���RK�MiT_�ʳ."Wc�x��8����U��7bm\�T�ܲ��N֩&�=�$�ބMd�0��e���Z�Ծ�p�
���4��~ڎ�)z���p�Q�5�@��e�+#k߿2N��W��I���?���� ��I.2����ӷԈ/���"���
�����v��������E3�����#:I|M��0p�V��`���pY����8��:���?�I��a
�n�B���<�^�����C�)��x�f%_v��I7�IEѯ~��ͦ6���U�wߒ��M��Q��������y�מq��R������;;��t=���vĲ!]:4$Oc���*6�Ƭڵb׍�e��\�ƜqBgk_*�
iEt$�D�}�w.�㧹�Ξv�4�K�6GxNTY	�УY*�B��@oê�
i>�,�8��ڷ�0'4���e<h_��H���մ�Ic�z�7�&�k��ê62i�������L6S7��7�'2���^-<沀7�cVP����> /_y�7���/�/���� Ȍo��iq�Q�O�Vʶ�ڢ�ool��7$N�p,�DRU�]���;e��� c�sy�3�EBK[2w1|[�����U'T�PZc���vo/x���f�*��@خ&2􈐢0X�8Z����1spU���|��`��x�^�0�7
�һ���NuN��h�SXsX�H�|8�H�N�vM�)Y\��-A�HJ��$/f�&��0��k*0���--%Ro�M�ys������ܚ;�_vD$h��"����Q4���6���"a�>��	9e����e�o�]4����s��%����ɦ���T{�T@T*�ל����+�i-��w@@#��R��J,���7����R�+�3�MR�]�@��B�*�#3� Ĝ�o�s�>�2,t.:�c,.h ��ЊU����h������ry�f��W���X2�M��>d����x���?�_<�R�g�i:�3��7�R����������kr�ԧ F/`t{w��9|�_Sw�c��{�>��L���Ϸ�qZqL7Ғڮ4W�~�#d�a�X�[�� ̀:�7�#�b�"�� �FT;��y���&i(#�}�>F/ӾsZ�Ҧ�&�|";[������:�T����oZ�F�?�TYz:�<���1��{0	Ϯ?2ep��U�H�Wڇ*u�(���> ��	�FA�˟o�e� �?B��|� �<vk6�6��M{�@�[9d�Y�׭~��ݢ�P��F�r�O�:&����aREl�s��E"����H��5և�v6�k�Y?6����9�L,U&=��غ0V
+���C�b��p��x�	=f	)�P2�6�r��4�C��D5%Â���`�0?�ϕN`�N��=3��q�q����5���tC�����<��ί�ۧeH�DM�"�H�@P7
�r7<�_�������A^µf�����&����-Y��<��:w��a��6�M��d؇!P��ك�\J&�l��o˞R(d���|��kG�_���_���a-���2	K/���􁁮��;ɰ����qІP9\��A:��ح�T��v�q�B|�i/���m V���Pŷμ.�9�'�ϧ��=�WCu[|۷7�t�j�y_���θ��
_M�ݕ�`[\l��3z3�֑76-j'b���j�Oe�BF��I�5�ivٞ�2�E�Vb��m�库�3h*@%��zP!�秆�� #���A�� �҅G����eטzM�Pl(X6J���4tǔ/��QoE$�+:)�`���t4 ��D����K�s=�JN�5���Zg,$%�7ʣ��x�7��a*W�A���܂P2߼^H��h��j���}�����f6� d���@��QV�'{�V��{ɐ��I�G����b�m�e�7����z� ~�ܿd+�1���Q%A�QA�aM�=���K�F�ٖ���^�/�>�U���)`�'��S�v5V�M���!�q`l"\"�0���m��J��\Z�ZE�B��31��6���@$K��Zi�c��Z����N��̸)�A�,��쏎�ö�"��ت�"q`DR�"�&8�Qܥ��@�b�i�T��4�O9&UW�Ļ5T�+Ć�Ϫf_|�<���V�L��Iع�
6�g݇�^S����O[ۋ�s��f��7�v���p��InE�/�Si����s16���|�8�r�d��N7�<��mzM1�>h=2���;�g����	`.�w��'�Ws�#^&�+��tPM��{
�3fq��LqU̖��m��A�-��GÜh����ʡ��`hr�P�,��4�
�t���\�$��{��+k�?1Dy�s1DE��Ceȝ�['�8(��g����C�鼼���m@�Y\֜�>l��s�/��JĶ	T��	�I�!_�.�%<ɛ~�T�|����$ks�j���o�0�}z�J��#�M71�gr��W�HU�,� ��~�3���?t�Ies��$�9�I�	���V��=V�����_��jE7��`�Rv�b` }�<0��e�:	�
xډ4%����%�����Zl�@����	�y���4�vo(D=�b
EX��u�㺈���ͅ�)���2�3�Fn5�d��YǗ�Y_�
w���]n8ft�[��z�ka�oY ��cm덶b!��6�lg�,r�ځ�XU��Y��h�ʚ7 ��������kS�ޫe�f�����tFG�9��	�C:Vߐ�"��u§�h�#6R9VA�mP9V�e�V�c�� �]����eOv�AG�P=R>�'��e�a!)�2BxC�ὣ
�Q�D��6���nPU��+�4�;7VP����PW�/A=�yy�!� �܊X�H�9�y
��a�����vE�� �8	qx���dʹ�EzǼ��0p,+���Jm�2Հ-�LT+�a�<�U�n���������:-�ML����L��E��ѻ\�NB�W!8M%���{U<B`q=�щ��=�N��q@V_?!�ۇ��q�e�~T���&���$40��&O+�E��1%�Y$3Hv�HAj�k�y��
�t��ʐ-� ��jlh@��WQq�Y��=I�_���("7���CE���1����i����[%�Dhnwf�qiæ��G�u=Q�2a��:	_̻���Dq'�ºI6����A~	n�W�۹�R'E�:��Υ�Y�p�ifQZ�(��-����RCXx�kv^zET�k�a�QW�ӊ�D��� �ڭd���8��R����`:72�D]K2�ܘMӣ���^R[���(�h�a��9�sl��g��o:W/�ܶe���0��a�5(��Kv8��mR��r��
����ә ���Ĝ��#�����ݲ1٭���4�� ��
�T����~Y1lG�=+̃vn�!�_���5Da�&�[!�@�-��^8�F� π�B�i��U����9j��F�D�		$�:-?0ʒ�Lt���aa�>1�����-6ĴӜz�'j�T~ }��f",�>���iK������!��1D7�#�s��J-X0� �7IGV���M~y��ՠ�!" �|{�����g2wu|>W0s��F�2T��[��]&����_�������-�,�>��ˁԂ{�����[�NR���[�!2�v�P8B��S�t�>%?"�y,X]�������{Q�'ت��´�"[�\�!��c}6���f�{���~Vߤ�4s�YiӹD^A����Z�e�������8�@/��8�iZ���0��HL����1�ȼL-��H�Z	��s.b;���z��z��:vu�C�57!A6�x!;9�'���&�*&bo/�z�������Es�����Eت�����~E-'X͆tYfل��W�]�QI`��`Ժ��y���jS�F��p��^��,��!"zb9��Ύc"w�S��._�@���IjN���Ju-h�F��|�2oy�%�d!�4T�cP�g�,[0IPK]�*�ŊH�MPlH��_�	���Ӻ��k�7�T�uU�-%Vɘ�fE�U��	�`�.�˙k:�㮮���U�:���z�آ�E7q`�8��Ω�p���.���{�t����Kg���g���=���*���:�!�Ȣ^12HY܆�C/c[�~n0��	��P���upp_"�5���D,�2S*+&{9- �˪�i n�X�D��Wh����F+�+,Z���}�Dd��_��m�y���.�k�[���m��X�H �Vj�嫋3�3R��S�R g}Z?��>�I7�2��ީ1�1�\���7�KI�߸_9��-�aw��5/��s���q�T�4b�������Vv�Ȍ[�1�Vy˿>b#�\]�P�k|������oR��)B�K�*c�琀l��옦Ƹ����s ���)���!pW����7�a�	(��#]:��ɵṁ�]�lȑ�G*1^;p�/6tf�j��+����r��G�ܬg4������%�E*i�X)�u�3M]-A>�"'����U�+{W�⑕�fQ��,�)t�"h�ι�Ω҃����e�e�B���1��zx4��1gv�X��8���m�>� S@q������a~���� ���74��M��j�щ���9)\kh{g�F�X �]�3L���~���Ӎ�Qo�h�t���ẕ&��*�����J��D�ӵ�2����4�����o!_7Q�/�l����E(x&w��N9v�� ��
�-��N��0��ƽ��EGE�����W�j��1���]g�ʺ�L}��:�,F�ζt	���hA��e�]�X0{
AR�R�@���ևm�(�����)�����fy���Bd�����ld�{�QT�R�#]�,(��-F�&S�H@����b.�O�"�Q5{j��L��?Ȼ^�.�g!ҏ�i���F���'���Q���JfW��֭��)1v_����n�Sݑ�[��|ha$��Rl�m$��
�k�qG�9��V>��6U��Jς��F��4�8ǖ�.]��j�����? ��S_����&�N삶d��0jq���C��L����i�s!��m��;��_�Z�zq7�2�[�ڗ���}3�;3�5�6�B���ɴ!��?Rd�ޥ��-��~!=����P�������fw�ۋP@B���s~��;a�RD;�I����\��n�+쬢�A?H�AԆ$�-�A�AO8�ꪢ���t|�����rʅ��_�吇U�����6�����J0��k��`P3�j7���-�_R�q@���o䇣��Y��rl���u���ߟTd��n5B"	��f���-5�qT�=-���d�B���黬�R�&���p���H)�R S���&Q�4��)���[�2&��D��A5u&�K�>Yk܀�P���A.�X�oHtjy��&�M �� 28:u�k�0���h*AX\���1k���kH�����Ϣ3҅��T�M�]i�2N�3Vu��ߨt�L��fS8�Q����/�{�8����,�}ԍ�Z5�Z��0���n9��K7�Z�*�2t�h�вǣi!�c��������KQ���KM|e�p9Y��i]u:&gV覷�5�\�)��x��Xb #����`|!��47V�"	v�y�E�������g:���O3��Db���ů�����^���ӄ^:�ab��\����3+!��1������Q��� 
'��ǀ;�̖�Ƹ����:Ar���%��\ԥˌ�Кۈ=ȏ��F��"Ă����-"{�?��8XXkۗ�':�C���>M���>�X�	z0&��h�k�b;rκJ��h�p������_aL.�0�Yo�`0����u�����;-Li��i��.��hN�t�k]�
����X|���i�<F�gH�^:�UDaf)�5��pw*T2B�u�0���;�t�:?igt���ZP2|�^1�H�����m�[w9���������IU`x'7�C��}j�
u΍V���=��G�j1���K�/N��@J���)~�w6=Bu+�",o��8�|����S)߁�S�	����!���>D3�}�3D+�}���8s�|f�
����w=�����$�5� �������+t��w:�0��t���~Y�t��TT�LeB����=qSEW�p���-|�ĸMZ�5��.ᏽ/c�[U;G$�`�o�d_V�!'D���4�eoR�*Z���	1A��fA��H%V�n�H����}	j�	��t>����I���=�q��D�l[�)-��B]R��� �K��S��n�^]9��;E�9���}<FZ����0���7�뙞f�T���1��v���[j�<#�WϚr����ߛ
�DS��sL�-А�\ȌR�7�\�m}�(Q�����'΁f3�k0�q�Ty1�7Z�\f��ɥ�La��A���Mi	��}�aB��ә�Vۏ�]� ���Ϧu�L���r�pW�	(�Z|aEr"�U�T��;kyz @�ߔ����B%h? ی&�<d'�Wծ�~C=Np3Ph�ϙ
�!̈́��,��Ie@9���֍h�T�[�������+�_�'JL��M��t�����9�y��k����IA��hc��{��Y���4q%"��"��a���!z�6<��8�!T�*44Um�V�.w��*/�0>�dW��ǲh�f���Fm�V��u�G�
Uh�e?8�]�_mt�U��޿.M���6>���Y߳�(�PB�n�|*�!����!ukZXr��~�|���4-��.+�%���֊O�n���!��#J*s���ङ�/�F�}�q�s]ԏ}�������R�YI��\h����GVn�oz�6$z�-�x�l?8}[W�1�0��}��!0
:�J�Y۹.#0}��*WC
Ͻm�����9Jv���6��Ó	{��X?�����˳1_3�1�);n����v��i�EB��L����9]���F��FW�R)=�̃W��^�g,|�\�&*���P�A�L�	S�}9Jc� �����x�A.K��A�����W�bv�`��z��!����I��p_!����/�	;?���=x/ʶ_J
m��wh�{~H�v��$1���z�o�J��-qK�
�S�� ߍ��5���1�v�J迩�p�8�baY+ot�1}*���8��+�#��kUs�a��:I�����c����YSmu���f}���rcqY1-Sr�G�����jK�V���%qHE� |n��$�.�]���n���ʔg��J\�����>�[�$A�,�����`"�0����/��:[�opn*ꘄO%��|N ���r)���)Z�)�;bWpj�j��Y�x�%��,4g��������-�H*̡O��?�/�G)}"a��z�@�nW�O;����S$��	�C�%����Dd
��LO9�4��_��;z�4+��	��A��]�uI]b� H׆r#�g¿K!�1���a�4V~�t��N��AQ?Pɀ���]�[4��þ��?��ҝ���Y��!i|�����8�����݂��7G@/n^a-7e'���Q�XDo�6�+|^?�²KIG4<�F�a�F��<�k�rr'��sY$V�Vv/I3'�ч��G��)�e|���� ?�/�JT!��<E��������z������d�ͱ�3�6Z�����|�yI��]9�#�Gʿۛ����:t�ټ�$���4ߚwb��((�<2응
1ۮ0�ҁ��+�(��M9���(��	�g���o׵�T�C�W��y�u(/��"� Jz%P�Xc�e���=�|!�O�fb,�r7���%�����jA�W(M��YPS�}�����Be����?:I�#?������X��<�U�� �I�#i��>�5|��ǝ�\��/)1��^߉eY�`c�U&�~-sSD�Z�����h���Y���n%G�}�a4�2�~��H�W�Tm�2{F�i�9l����b�}e�l@�b�����qՏ},p�� �r2��AX�a����gF?:�yߕ����4���W�6)�+�"�\�_���5���kF (��I��7�|�!2q9��z�q�H�"������ܠњTcG�G*� 7;+DXl�[}r��7�kH�@{��<Ƨ�^�jUs� "�@�p��c�� ��X�<��%=7,�a�7ߑ�c��SЎ��aod�QO��2�J�Vlu��N�p�^
�<�c,iR�j��P�u�v��j$�ײԻog���V_
*$��H:u�@ݦ�t���PF9�~j]�}��Gf�``��7��H������u��{�Jl��ws��&[	vh�2�ww]bx����g�'��\]|DM�Ɵ�a�t�Ϛ�D\H�عۦ�'C���d6�x�RX���yae	qBk��$soM��!��oM��K�0�)�r����t�|T�����rR�����8S�ի�g56;FQ���W=��i���
�є��>Ϗ�,n� �<���d�D��a��0��̑p���c��8㯟a�9�-�pu��W�	�ó������y�`K��|%Os��V�2�V��1��H��S����#������ls�⡅B)��K�/��^J��4@.'2�ao5���B���C�����	�n�F�/�]�J푾�?hP�_f#��oo/G��,O
o���]�O����lVc�a��v�S@俓��PJ*=Ry_�.��l��l���"�g��l���8�a�~v�p��p!f�Yl+Pl/~��_�޲�_f�>%7��.`d�z�b��/��[��Cdi�P�
��?ޜ��a�q��>_u�E{'X�o�uw�+�ȼ$��n �d�'�es?�A���B�T�eqn6M��Vv`�]��"ژg.�u �͙���c��n�I���)��N��F����pc���5�%�J�r��3�H]�ǫ�)���[W���԰7Y��W'z����Y%*��QVV�}�6Al)�����B�]9Z��%�G ��	������������\N�*�4����)㾁���$6����qI��E�3q���;<Y�����7K�*�'	���3�����8~�tA�!ÖG���grvM�N�@��l�L,'i�'b�@9���M>� F�/������u�4���>�-��u��:!�V���Y˔�	C^I5-��1�m��
���\�	U��U�9W�Ahx�-I��C
x���i�s���Ç�E�"`�`j�,*,ϓH)�c�������RW^��˕�!��n\H�5�����e���H<���Q��VpE�j��_��n��ʀ�l�X~S3s2��� �<ٽiT��9W��H%|��ʹ��oӒ�Rq~ �7��J��M'��F;bՆu�%��M*1ʝK�_�aJ�[�-a�ѭ�}9	Oç�'�O;P̡U��ƽm�f#�ݙ�G��z�vү��o��I�E7Ŋ��t{/U�ڀT,�V/:�K�kR)����-��{�8|��4y��^�N�m���+�6?WQ�LR�k��މ�O�����j��GŖ��^�P�W�R'�6�W� v�3����qR��P�إ3��p`x���j����ϒ�etV�Os>�&O���YO�EJJ͌9�I�P"@���%�=Kq�}��~^�ƈ�M�5\���I	!�G/�н^vK�ͷSo�s*m��9$�UY$ࡓ�fGU�E�J�{O�e	��G1�K�{�Z1��p���U��pud]�Y��tUkn1@�P'�8"�q�|V?4�~�W��=��E�CB���]�/�HK7��sA7Z@:z��?Xx��<K�:��433(G�I���*��d�-��2�b�ۢ햵y# VX+��2�X��6����6�rq�N�����' �[�ѧ(��ݞ=�c��88�i�!�[�����Z ��(�P[$̩֒�I�n?��L��OB��"�h�Z,���c�U��I��.3s�c���h�1��K%�H��L����+�P�<x����QiJ}q�<�ƊDyɂk�6!�~a_pj�K?f���+=�ز[nٻ#lb�.�S	򵒭��g�
GڴO�[�)��A�>���<C��c��KBA��T^_ӱ���[֌�9�8)nA+<gn%FU~8;`RuD����4>�na���$�C���oܹ����/����$�L��������y�]7��Mŀ����^�-<Ɏ��/�x=��s)o�=}��ీLq�����0�|�~�����6.kD�y�m>�̍���O�(�Uˇڄ
�� 8'�~��/j"�\
v�e@�E�͢,�����<i𜸯S�؞g�\y:�f��8]K�Gl���1�%�x7o�h�,5Y ��Ӹ�=�Nt1V��,��%�oK��	�DCwF*�t�g����z�As�0P/�D5�gr긯�N��ݶ)1��vAi"{Sl7F~�s���Y)���?io�4C�9��4��l��!�%T� �W������m"�aUH��O<1��f��_[3:��>e�<Θ?�BE�{ߠ7�Bu��Ǖ�H�� B"Uq�yW���FE�c  ��q�p�f�E�@�Z�li�� �P '[jX�UF6N����.���}3�c�3����&Fsyx-M�E`+������G/��iI�>�f�g�NӦ���*�S�	b���c�fN�9�m7s��1��}^�P���,�?~����,����u��9�� i2��
������Ǿ��<)0L��nlߚ�~	T�H�����èt"�L�k̤f��j7�j7�V"�eC5I�����B�Ġ����������A��p"��a㢑EX�}!���]�E�d�g���S���ǖ����j`5x��B�b�¢�& ���ې�b|����!>ә�� ��Ϲ�ΰg�BO(R�_t�~���j|����f�%�I��i���?g����d����n�z�ZeQ�@A��\M0��1��۟��so��y;��V�%��������xx���`����8i��z,%�E�"�������Q��^�N���XCp%�_�D&`8ܞ)����|'#�ۛ˃�%R�%}�=dR0��̑�<��WX\`�ݕGh�8�H�k����	s��NɃ��M�����Du�#91�r�EA��֙�X�nP��o�qTވ�����S�l�*q��1�?�[�lU�`��RD6,����S��YRX�#�W;.��s.i֤����1Y��^G͜�p ����T�8�s\��H�3Ⴧ[M�L:��;�E�i��L�ϓY��d�"�/�aD:41%@i��V��
�A5
�K%�0ᖈ��(١���Ƭ��V_eG����/��(�*k,St�d3 �� -��5L��ʑA�X^�0�� *���2���n?̘��;I�r2ˋ9���2ꌷ_��Ox�XS�vD05��PNV׾��+դb7mL�gR��ąѨ��9}L����"���}��yBf��}ߣ��*?4��:�f�)��r$�[�	9�"�^��1~C��CR��@�Ƃ����76I�:U?5b8d��_��������sޤ9���4��_�����{��]���`��B����Q��Ԛ��Ei|�[�p��� ���>����&9�~_T�2��K�w��͏�?x~^�����l�,}��m
ZC&z����[���
�7K���s���A>���u���y�$gX�`�@��(�vFM�4E�ɧW��>D��n �I���G�!v�,Şъ
�A�I�x�ޥ����ո�O���/�oJ�ִ}v�5��4�%	qg����$��n5�}Ɛ�㯾9���� ���:d��@� ����^R۴��O%��p���s��Iy��TA�AN�˔��s��6����W��l��#���
`9�fYX��!ֶZd�2"��-����V���¥y颼���]�T7��rF{h��lF�!,TP{9�ó�uma�q# �RUL�nR�v�1���Է�Q 3�\lX��������2�� ��,�խ⮷a�Dzn���ĀpU ���!����NQ	?es14i�@��\��.,P���)�p��\Cv����JlL��n1qET*0�tK�(���Q)��S����y�H��Q�Ϲ�V����*D�&7W}�6͈�ٞiô�,�t��w��!�d��#}5���f��j��<���F�~��`�=r�n(�{|������Zw�Z��2^�܀$\$ʇ��]���<��oo�͌ ��2��A���n�������S��oR�x�ˡp�F��e�N��s��)���^��{��4��F��7��e#n� �ANQ��s9�L��j@�>���^3m ���/b1yc0��]`(��8y9��x�[���rq�?@XP{V�t^�Lb���o�^��&A�a�&�Y1^.	ߗ`8fS�/%�&�RT����%j�����W1���E�W����	�������(�]�I[iJ~�9G4UsO����E؀��}�s�r�="�w�¥��w�(6��(���F8�"QJL�~��ƛz��|?�Ț"�Hշ�M��݃�W�!FNY�[�w�d�.�;����q��B�Y�����`?��g8uϮ��k3�cO�4�*�� )���0��9+��'v4]�v��9��@�B_&E �'Y�k�r�G�wd}fz=�����6j��j'=ʨm����D>�G������s�^>H�?H~]�Kf7�8��+h�d���Jk�N� 5�%m�5������  ͩЏv�yI�`���U���J���N���+��ڰAM��v���Un��cǦF)>dḒ/'96�?��sB�3�S�؆3�9<�{^Ku����Px{��MQ2Ө���T��۳�O������7��0򋠊�T�OT�3u�kYѠ��u��6;���t��c67��T�ǵ�cѠ��⌹�����2\]Em.؀��$o�Љ)U�N���iM��I�(ߗkP���RC�Lm�tTdϘ�?����bҨ8աƸ�Q�&k�	��;2,��|N��H�|][�Ik.�m���1Q��}U����<�b�����f��IO�Y��А�,�a����6�_$�&M�iȗN��U�x�ƅ8���PX����*|X��'N6T_���ӏjvU�$�����Rִ�yl/�	���H��Z(�(
�V���,h&*�Z��ԛ_j>pl��Dʳ�����o�f�N\�����R�S�1���	7#��n�"z�E�pj���U�[f�,YsJ��T1cst���c��G���A(4�iN��|��Oz����1���D������U��^��<��B���^P����t �z	�M\fz	�u�\)�����[hh�F؉F������tK�m]";�����L������Q\�p�j��;|lb4Y�� ���V�����<;�]}��|S��h�"|j1���ǹr+�N�_�.�o��X�����ٰ��&G@��Y�:hqV$�aT�u@1��m�T��r������oJo�B���P�$���/���(ݽ0}lJ x	�\������9Qچ���,�D^��k�FA2ړ�F=�����Z��a�!� ���ҏ���f(����
�2��1�_B9�ۃ�TM�V��*{��H�l�p���|,!�-�7-�E��O	�t���Z#�S��Ť.-Ӭ��i�"��ӟ5xB!�'�D�͌ �$�CX�`��u�K�-�D+^�gI^|Oa�&�ۆ1���4fM������dJ�я8Sr;���/����*t�yD0���}lU��=�2�5o���z�Q�v�ݸ��/��W���vB�n{��B ��m%�� ��σ��EȚ�Z��?�3"T(��A	��zL�m /�S�۰S�`�|�|
$�VĐ�t�p��$_il#U�Xm{�Vd&p6�jj؀��*F�UV�h�1��"����
PF����� ��>ꕩ���l0���Y?�-Ədv���-O���&z�����{��6�{�Q��N�
���La�0j�.�A��ª�Y�"��Q�HT��=���E�Q|}~�$��/歺�s4�m۩�>�>q/2�m4�ӳ�7��T��ql��v�袋V�z�5�>yl��ж"^��YB@����-ƀ��n��8�� J�`��6�8NU*�+��oҵG��VP�Z���?>��pk4�����:�����,�ۖ2lS�.Ċ�F��B�����q�b5w�v#���I�"�F�[����ς�R*%��nI����Pq��d!J�tQٸ�q�:Èו�?�d~~I�@6�V����$N5�oy7-���{�O0hs�
�(��鵢�(����l�n|5;��e�CJDՒ�j���|��ƹ����>x�Jà��g%ǉ�4p�w՚5�v6�e~>��r�J�/�,@9fy����X�{�ל}W��(���OIE�xe{�U����{����n�r2��՚<��F�������;.�?^,�<D(��6�ޟ%��琢-��-���t�ς)d����S��Y��'rz9��J
���q}���yY��PG�p7q	;�������ƴ}��o��E�v�����5p�;�Q!���O�Ɣ`
�뮇�|r�4Θj_��=y����3��F�u���s��.E�.֕ I�?������������K��ܗa�� �����'��A>Z��F75
�4ˁ�8cw&�q"'eʰ��T�x�ôASu�5
QH,�q{&waۻ�}���:��Z���.7 ��9�����@��	�N,�����'�
�x:#�	����t�����{��fP�dN�%�AB>�t�s&�xJ��^��*w���?�J�p��3���9�aܢ��ⲣ]�@hqx7� >����FW���:3�+u��\�/+޼�r���!�;��O��3�� ��K����$�A~�FK2�l��e��
vnejg!�x픁jX����He�B��	:7��y��eȉ�dy	��A�k����&Q��K�4�50�����PB�h�eҬ[G="�rɜ���F'�f��Vy��N#��s蜨<�O�5���C|�b�c�x/���C��=E��Š�o���M��ݺ��8U:n
6�S����%	ЅL�Y�tH3a�����}�C�_��*�G(�M/fk�HR��Y��Kb ��3Q��	���|�5��s���qgn�]"0p%�F(�a�;@⇫6V����K���P��d���@h.��bب�,t��^:[��D�މ���M'�cb���<�pggl����f�.elͭ�n���k���z��У��`��@��k��~��=�Q�Ud���n���A���a��<u�D	����f,�xK�F���R��j���J�B �Hn��S�"k��Y�Πqqب�P��Z*LG����E�hW�\@ʽWۍ�]Z�,n�2�Ul�=���QƜj~�E���E밉�s�)4��π���E��c�3e�nR,��^)�I;"��4ln�����Lo����2 ��'A�1
�X�����~����ւq"r�Ώ؇ʹh ��\Z4:��,S���w�	��m\qwf^Gwq��s[bg�B}�ۚK���^\-�裈�ؾ|��6#�c���1{cf�2�G��튢yWF��7j�������h����E�-�A�y�Jpĕ-���R@eƫ��v-�����H�gm�o�KU�&0ü�?O|0��/"}��R�
_+w�����VM�^�l
st�|��4��\��������`��z랩ւr���o�y���^��#Y)�"��:[��W���\E\7F��w�O�He����j��qO*#�����F}T=9�鎣���&�����AD֌�.��
:�Kс"Icy����	��UR Ɨ���v#ڒg`�A�W�sb7��6�(ի-�G��9�����C�e-v�L��]�%�1�(p5��O�S]ַe6b���R�I����qI����[`	�����L���ɽ�!>w�����^�:-<SA3��rrhu��!�����]�ǯ�};����H֔�T��~鞼so0�����%q��ժa.��["�Ss�OF���kHR���"��4���3�p��3L`˵��i��E�wlq��E�)~��xIFA��""�])R���AF;��̋W2BU ��tP@p�U�N�#�3մ͈/��X���i �K�O*r6��	���7\�zzf��*�^F�C����c��2��IkI^>╜<�G,��gvh�eh?��3�T'\�%<蝨_.�0WXD��~bj�������z�)�'�
"��H�p�{�!��d-�0��w5�@}n�AIh��~해�
�g��m�R7���l�E�A�%W�d@\!�N�O	e ;�1�R�/b�8Ze\�#/ ����A	z6l��f8[�) H�k��9�w��������r�J�\1���D�m�d�N�J:%%���)�y�U�HmsDq�"r';k��	�l�Ƅ�NR�-e�B�p�Zw�8�B��<��+�V��w[C��%i���]�V��uuk�G�6H�K伩�	W6v�7�g�:�~k�����"Vp���&�S��!�e��>���(h�pN��ŎJq�/pH�h�w^�I�1�'=���
:E]����Z����iX��{~����2�s��V��y�O8��Z�e�B*n�UPřYLq9�:q�)`�����e`��2f}���Z��Q#�7��m��єF���8�yb�[=�K&b
 ��'(4P�]���B�%-ի��-W"��_�C�Y��{���괛�t�5c'Fq���Y6��/w�!�m5!϶~�R/������|���gBoǾ����`"�d�Q��S�1���N��r�̒W�)S�vX��Nݡ�\�@`~-&�c�b��ky&�I���*���Sf2jZ��$C#�B�r�������n�PL��.]�1�X�T.$�,����JeG=򌗀��+�a^����P����2?�m���A��6�3�8��H�#��L�+Ǽq���*�� �����6FД�|XT���k��r+S�8M�z��
>�7�"�����U/a�V~�aV�үLIv����jRǔ�V�����t_^��pn��Sh��\�*�k�O�`0�k~8z�����#1�{�s�����!k�@�M�Q@�#���P�n�M{�
�wtM���Q��L�'j�x��Z�H�l��C�a"�9='��Ґ$Fo�H.Tcp�b*�P=���ב//������iRFa1���l�c�A4hOl��d~�<�X���X�n��PJ��!��$<����ϝe<\��mT9� i��u��]s#l�p�1�G��k$b�52,��z^KŤL�	��~��b�g���a_&��9��>�"��
�E�WW��ި%��P�z�[sS��z��i1_Ro�C�wP o�N�:0�|�3D��I*4/d�X��٫"�	�t��O㪰
�T��KHf��HQ��｛s(-�9�L�(�Z|1�s1�ׄ���9�t�@�CI ��x��&��]c�$��e\! ���ۗ�����O������]֜x*�貀Bl���,m/˔��8� bx~�qK�h����s�1�*XE��/�pU�Y]+ro[=Mwj�9b?%[K��qk���P�f�w��?k����uq�,�Ď17�T�Hq����3rdJn��z)3��;����T��0�#$��<�d&�;"��V�;6�o�ꖇl�C�P^ӟ�?������+b�cx	��w�2�)"¥Q��MS����(�k`���V�[�×�n��|X�`u����c=�\g�&d��Q�ͳ/�)tCEq��GsPM��4�6`x�UJG�ZFv��)�Q��z�����A60Im���	X��;����A�����vޝu�Уz���z�� �a+(=+KoP7�~�ء&���'�pFU����\�d�5!�m,�W.�+��v�K��+�Q��q[Pw{k��Oԫs��mV��Q�OW�)^���W�֡�� �,�Hh��0�1l���uBp������?1�a~H�q57.~�辘�E�7�{�_�*0o^�JYt� �V>lY�j(K1e� �U߼�7ʮ�Fk�Mٌ��	=������iZs�� � ��(�Ȼ��h�K&TN�,���(
��+�>I>ru�YR^�y�J��K�@�y29Q�bW����yH�@L`wa�(���Ě�\}��nv{_���Oq"��U����IO�4Z���M1Hq�BN�u[Hs^���2c����+B��&Ϭ�9��62���l)z�K����o� �:a��T� $�V��,��&��_��|,��,}�d�sn\��@^�н���G��͊O�o�j�p�����C))Ѱފc�<uƜ0 -����6Q,�Q�h*���.l�b[��#[͂�Y_8��zȻ����I?%�L�C�RIP�ʙ���|�
�I�w��C��u��hM-S۲o��vMN}�B�7���z��f�M�臈 �@�_,ҟ��Uʼ	�����%���]��1$�U�K"��#̓�X��xd���t�]��|߁���=�����8����JH�5T��1;���JDeR!C�m�fف�tv�W>�h~y��;�ŧ�?�2|4����djX�N��w�x���%�b���˓��<��o�o�a`��#�s�m)�1C/��9P���0{�������.II�/�u.�H��*f������;��Ř�,9�A�f`hZGGC&��ǀ��Np��X����ʊ~mH$����g�Df�*�a� �q��c��@�u,�N�޵��78�~�L���ť�q�=����V�vV��^��$
����k@Y� xiO����ː
����VaK8ps�~��8�����e/������Fd�FVi?v'�.�d#4�?;j���Q��xj�T�z�,cP09�Z�&,O���a�c����{T��K���-q�0������x��B���t���(��KdqH���@�u����@��p��>��`:��(̄�u��VQ
�w�(1#�*b-�:
O�����S�Sa]�pL+ʃ݀%.�U䗵;jI��d]T�Y�U�H�\���E�E��Le^H	����wxÂ���
n �ݾ�Ґ�P���$���͏21V&�\$���6�O6��I�sH�̎�he�a���9L9�+����.�Y/��}1���[��QU`�Mp�9���vx��������R�t�~F?��pg	r���-MÔV�eos�y�MU���E~M��/ap'=K���!����gq���3��y�ppWK����Y��:3чr�e�6��w6�~�*E���b���*�*��;�Q{K�S��]�}�eL�&��-�ۏ�5Ӄ�����i��s�%�c�>xÍ�?b���X.��퇖�0��PsKH�`�w��BMo��DE��-�"��"�U�̫�p��O�w�� |h�@-���'��.j�O��BI6ŶF�򦐵9z� ��DR��by¼j��_����������l�9��R�u������@�W�;��E���D9�\��y�����)O��Ȑ�Ӷ��蜂п��ʲ��L˰�M�S@�l�����:�H���Q��Y���-����DJ�υ�;Z����d�`0�f�����D�$� ��j*,���n�m��V����{�)���p��^���J�sl�s5�q�{B-Z7����4���Ew�u���� ���AN��o,�lZ�a����%c���1+1}ú��-��R)p�2�όN
}��J�/ط���l��N���Z�yCӉT�lh�k�S�l1�S�h������0�B��c^j��厕O������V�r�l�6���1[�H���Ram�Z-��=~�^��Lq;����ASn��ԥ۱�f��l�w^h�K�x��s�I��H�on�&���_�?�Q���BN�A���Lkن3�J˅d`�-�[^1`|ڰ���,�Q�pb�=
z�s[$ר^�y���/|�_���$�	��G�8�iYEI����X�Mgx�P'�~�g�%+�BYcc}�fhp�;PpoO.3�K>��\z�ȷ�|�v��������lM�S7])������:M�-�`"������p���j����`��`R��[��<�Ni��k3�`�������p!3{Ws����A�g1�
̠�L+��.9ñ;{#a�_h��m�穈��\2�FL�B���k����D��TȠ����oY`��[1z$��q�v�x�׵r��
@�
	����
I�Uf4��4�2:����a�e���D�����X�8�x�h���U�YM��,�2!�x<3.(Ҡ�LLuqG��!�W>�9�.����YwT�r|t��7��;� �j��h��bY��V
r��QW	,]��M�i��1_2�M����T����Z��{kC^�{gc�r!v�H�L�3=��i;KLV��ң�9Ҭ��������<�����V_b�.�g��A`�b�Ʈ���\qk0j|����!Л��8�n���ᶡe�Y������D�if��[�%��Ra��� Qt����0~�R���zg9h�X��@U�Ə�����.^���V�c!�ì�84^g,��
T�z��s��F��AV�n ��1։�D�aaQ�: �p ��x!���pEN�pB ��Ψ6����̩Tϯ1�X�>�hۮp��u�]|)��~�X\��(��ƪI�iavUO�7���T��rZ�:�am�Om�-�)�fbA��&��/4�$�;�x�VԒ���[�oO��*�9q9�-
��m�7����>���C6$YG3�B�غ3󖿆�yvEB��f}��Z�?x�[�a�a�T3�X���%�����iZd���.W��e%�+��"���(}^�K���'W����\���ƀH[���
ͺC�(����5Īc�;x�Msk�Px��� �Q�Լ�_$mQ������FM�w0�O��q���ǫ-�����[e�(j.��à�h��~��/��wb]�D����եq����t��Xt�7��كD�!�M�K��w?�X:�#�!����~^�����[�ԂL�K��5HE��1����n������!��Pԝ>�w�_�hG9Τ��x7U�\C��t���
� ],+�b ̸X�א���?+��.���(��Fm��� R�~d�Q�٪�og����?ouM��[(31 hY+=�C9�<�!"��̣d<�O{�>���5�+�
�����X��)�&ض=��x�ue*ݭ4g;�~'�̘�_ǝo�u^F���w��
	Ư}$��e�pzW�G�a3"��vV�i�\|9+�1�;�є�sma�D�Ի5!�vN���Qp*},h���&���v��7�>(��sVo����ʝ⇶;4�@�F�M�,?怈�<�=�b91J�	Γ$L�d0�1w�yʟr�u�g���*���:�XK��d�f�c95�� Zi��d���Ї�1@)E���5{qL�0��;k�������9D"H�[˰�>j���E3$�65kܭ <!"9����LJ�ȵ�=���	�~�	E~�Ψ�e|��ִ4��a��	����zUZ�{颢8����x@	N�R ����J����B2�O脠��%�
/��8�Ǧ+5�iTz��
�ժ]��#�u�4�/��@�f"�k}��2P.��0J[{��w�C�a+d �X�@��y��R�ߗ̒jwRjP��ϭfP�O
]�����������=đ�[�D���N(.~��Ǻ��t���+��U�%�А�.�]���%K����]Q��sK����`��C�Iۘ�]��PC�s�s�c 3y����7���7t^Z'��Fn�
�>!��6k��GRZ/��<��� +�E�����ٵl�+��p3F��a�l��Z�2(����H���S�R����s���ҹj�r`�����'�����u�_RsHa��Ϫ��%QN;�~����4��I!��,�o�6��Nkc���L��#���ך��D�����`Q�g��	l�q��H�����Wf+��墋���2���o��D,�|S�;]yn1Ұ����8{[���
�o<s��A����	����j���N�huJ�Uu�sչiCp�ݷ��	+o���T-2�$#^�iY��K;T=G�����K�NY������A;����BL�m�W�xb6%W�"ˌ��!�<B B0t����M���Yg��M��&��H�!S�<gF/2�O�(��4�j�A�=R�qV��$�^��H���]D	��9E�B@!��	V���hwX��tr����#J�����tD��{��=J.V��{��Ҥ���p 1q�@���~��I��ۦ?wbj���G�:��˱���ժ+�x�#���w��v�)�T�� tc�������e�13q:��ٰ�ǵY����Qm�F_�`���,��SЂ)�a
Aؤ��9�L�8��kW�M�r�ʕhUxv1`�0V���yU�ʖ��1��]�Q!L��X��]Ff�Vr$UU�A�w#�-~Ӥ %�!� ��y��<��`�x�������E�a_���9��3
-�Š$	�;;Xʵ�敡�(Z^���* ��X�vE��Vw��f�A:�P�z!�]#�±t%�v�{�s��w)-�٩?M��5ٍch<Z-�3eṾw�VA�/�U��3�.O4o`�f��m	al����w�/�x�hhk����s� 0؀Sކ��M�o����־�w�Q|	%��]��0����if�J��4���%���RB(�F���4��!�5�?A6;d��� ����&�z�����`�" g�;��N@T�)�]��0.����O����]�jݯ�ƶc�&ѦOa��֠����GTMN8��e���҂�Ĳڭ��=[Ua�������tS�4�Ώ���3�[D��zBC�����ɂ#�d=4�?���Ƒl�eЖ+��H�ZYF`��E;�l���-�������#
���#�s����attL�v���9Q���u�� ��\����7	\����IKdf�~���j�W<d��B ��Y�*j�as��_�ī*T]����|�[F<qKEp?�@�����w�p���/~q�����'����i��kɂ@�b�&Ckd\i�l9��TP�)8K7��f\�b��8�H>�M#���������_Kz�����P�h� �c�,����*1f�咱��֩2Q�R91��w�,>pL�c������6���G>��,5�Ɯ~"�1�ɡ+���t�|b�M�@��چClCQ�3	��u$-�à�2�ӕ-�=�Z(�n��ԃ����;d�s��>�d�-��*3	��FQ7���r�فK�<�f��ꦍы.��$v��]Tc�1=Y�C��:�[��p<����t^������-Wi�[%M�
/)�6�3v�AߧTMT��K�t+'�;�3�9�9�`�N��b��M|��|@Ԅ��������^��F�������ﶖ���-��G:\�^��m�n��,�3���b&p
S���h���\����H��D��g\ћ�m�� �t��A���/��٪�ˌz]]�9H��ADY2���;5��I�d �>�'����%�X7ف�0  �Ӧ:[�Q�p�n���@nOBj��)������k�$��2h�Y"�S7���\}^�3J�a<��F�����m��b�1D�<�S���Gd�}o(J�S4���T���-�]�j��ɳ �\���3BS?��Bes���y�ɹj$���^!��#*rS�@lCp+��Y��Va�U!�$�9��� v�<:a�����B��R(�Ã���h������7�1�%���HEi�B277�*3z��� �:����M@l�D6�ᅒ"�8$�n�2���ʇ���@l��s����V���Y?!Ha�=� �R�mϏ�j�+[ZM��S�]ɵ��j�FG|�	��{����7��:�:����$��p9g�ay2LzG��*#��/�7ihO�����BS���}"��ƽl9����1�4ǳlޅ>խ�me]16�zFG�Ba�qAe��\��Yj�'��Y�P�B����hI�,J��[�?�ֻ�~���/�����#
�d_'V�4k�؞�� L��k�'��s���*Z��^����q���֛]�{��P�#@�P�bI�`��Ӕӭ�)d�����}5T-��4ӾCM0q=�j�J�3K�6��$�1�W�񖿝I�EGBC�:3� �A6눧�� �1o_��Ŧ�prn4C�l;�ƀNW;����Ej#S�n^2{m��0�)O�d��L3J�0�r4~�A=����8F\������f�"N]�۴<<*ZCb�p!DLK,����U�ߕfBb���r�����:Ġ����]�>.���~ӫ�c"��
/�fS��R�%sz�'��w��q1{����d��D"G1���;�2���
�M^S`����)�^U\�_�[Dbl�|��G1sW�q����l�V�kN1V��� �ב�����þeLU/���k4��~�ޯX��#�}��s����\�/-i��i8^P����:Ѝ��L�}����\QX��}��dY�<B�`�Ǣ.F/^s&.��l5-�Կ����+���JF�ir��'iI�>�NfՆE�}N�E@��f��u����$qAv�4�Nl�S,�x�=�m�h�~�&��2I�I ��k�ӽ�.���^�$*l��� 3�K���da���'�����\Y'e��(D�
S�"��� 8��I%]7���`��r�]l��dUtJ\t[B� �:�1�Ϸ�hS�X��9��(��E�r�g�W ��G����=�z ����q��Czk�Y�}�� |A�E=�(��2�G�K��N?YԽ�*௧����F��$\��l��1X4���h[J}�ŕ0Ҕ(^�2���G��3�)��x^��ԇL'�餏 �e�fE�<���O���5�?��)�Q�?ɗ��z��ʒ��X d���yM�:�$1����	�������GPɍo�}U�(����dZ0�j�uJU���@x^��z2�ͻ�/��+�a�K�@;'\�+6�}9��+�OF3u���J�g�7TMY�a/7�:h?�/�tH!*j������K�I��#��j��Av�v������,o�%�HF���(6��bA���q�A�����t����ťh��\#�r�������[�82�50�"yo(���S�v�n��75/Ld޾Ѿ[�
}eAJ}`념�0�$�X�ϻ�� ����+��%P�Vݦ�rBg������LuK{�c�z	`��]x�J��׻��sуP7����ތ��h,��*�il��@� �PO���%���e�b����ACM�Z�%[ҙ
	</Z�Dx�^*��ڛ�L�BB������Mp��
�ic�E]̢�}������=�Y`��;�NG�'!9�1�������Z���LF=+���kp8X��
6����1^=&�n�Zk�3�y���x/���~���`���c`�nvx2�9`��(��8�*����u"�]�� i���' 鋮s�s]xD�J�b�A��_�W��^�����k�Hٝ	�o���N�%����;I�P7��O�����zY>�E0������҄�)�݌6{�Փ�E�����3\�v���7��,{�2���{��E�Q:h��WRӹh��/t�:8W���ӄ�('/M V�B�y2�w׉�;O���|���d&�v�,��M<���+c���N5m����s�X�7�H'���o�s��P92h�bf_��hĜ�VS~4p���\��d���˻�a��)�ݲk�9�0yhLՉR��br/R������ ��.�iw�A��\�S8(@�G�:t��ɭ����,J<�����:ዃl�QZ�!�wN�n����S�6�q��1 9�w��[�>�b�#,���X`��-vw�s�R޿�T]�̍d¬�Gc��&c���[R
n�Vt�fr�f4���YZ��*F�k#��Z�e�0I��CL�:���U�vU�i�"�����Hk.xC�S��5
�5#��X��AC��<< �d�9��H#�ce���Wv�wOD3AQ���"T����[�ň{C��'��vֳ�m$7��
c+GJ�i�G���}e����ܼ�gv:��<�Y��������$l���m�|d��|iV���!؏P)	�0��5I��ܰq�u�ln����@�L�1�W��3�Ar 9B��՝��s�	�� �+�e�X
S�;��	��9�VD?l#��]������(ʮVEx�]�/��k�-�
i^7��JP&A��7��o�,�3h��Z*�(ĉ3 �Egݔ��>fa�I���\���  e��#z�?�7D�@U�=d��ۅl�R$H {&Ɨ'僴V|����6��	ԲJC${.ł(!�_�坆/|z�,�_�.��Rh�)�J����u�O!2ʕ�4�R&��ޘt�h�H��� ܖMR����T���-
m�K��QI�6�v � o��<"cU?�O~��b��vV���`���Rӕ�`���$�G_'�M��3 �o�RkD1��V �5~�ҫu�5s���3&~%h=i'���5i���\
-�kQLc��}�,&���y��FKI�r	�=���s(�9(����� H���kYڭ8vk���3:?:|ef�*P;�BE���M@G�I<|7AC{2y�� J;�9'��D�)��g��(������d��[�D�N<W��*�K��m��RSΜO�w�;v�@��(��h�x�*_!�ɛ�0��aJ�+��>�ZS��g�ޟC
?�w%;�ak����}����GJ�Yh���vvӘ�f[�65cD���>�]�ݽS��]vh���n�:��1�ِ6�p�$A�)�aAB\|E�7�}���� 0���!&!�l��<B�vG]� �6'��Өm���tű���
���L��Z��QJ�(crq��g��U�S�5'ڦ�T��j����y��5�������37�@9�;Q׾<�،����צ�D\���|;.����H��˝�N}[L�.7��H���o-ĤY�����u�c{�ɣ��C�����(�6L���1	)��9CFE��}Ϲ�s��U͓cf抐7х9��|���of�2�����) -���`�~�5g�9���EΪ�	leӳ����T�Ǒ!ь�|�͜��X��{5Q`���S����u�v�]#[�����N$�e<?%FһX���d��x�ݻp8�}�j����=c�@�~��+����xP��y�o�Q��o�@����J��������ݣ�n#�g��xmU���`���Rɘ�xf����g��hX-f5���ሉK�A�ǎ�U�$O_��M^c�*XZI�$b�N��؉����2 ;]��]��a;�p~`��!�}B&> ���Kp������!���'�*h�� ��#r)*I+H�͹�� ��m:Gc#�G'��0�b�!�� nE�L��c�f��3j��Q����)����q}��C��w��n�Xٹ@�Á���Z{�h�93</.^��Ǔ8�Y���n�NNLT:I�Zm��$��Ү��5�r{��r_�%�8��l�8dQ��oG�����h�+^��qH����5�i���Zl�b����){-���L٨T�;O���"�4�`�-rP�袦��DLި�<���!}|��Γ]b���5T_�7��m��6��c�����fl�s����_Sw<�X���pZl_Ͷ����:������碮������������� mC�vv�kմ��*���l����*�u6��֞�>!9�4�*&��A�Q{�Ӄ��}Y����Z��M�h|�+/�ɴ�=�>��Uy��jd:�'b���{�T�Ѽ;5����ڧE��Ƌ�(�K �L���R�R���d�9��J|��yA�)�G��,��~�_���(?�?���������b@ �F�ɡ|��-3�up��E�`¯�W#��1���Jhw�� �9E-�a���iw����Q�7����xN3O��ƃɇ��r���ːp�q��d�}@hVC1����P9gh�o}�}�{,"�(;��6_4������p��(�H�[6��M�$�
����]������k�x��|��	a�sI����PKzL-���H�L��ꮢ03��R;y߈�S��	�%c\�A��=cH^���:I�7��P�t]�
j�>C��;ݫ��(�{�F�E�����#�H��H3�UKn*��ҿ��E&��}��(W$��;��"��Z>�Y u
��~4�!�������-Y���ɴ*E����� ��^�o/0�'sG���Y�d[O���A�<��5BTGl��akHG��xZ�B�2��"�p��Jw�
|
6_v8e ���j�־ �3_�v<���� ��f7X�m�]9�d���ѦNw��p>������q��!K�)��ןt�JdM����'�IE+2u�}E���p�����k�]��]�O�5����q���MF��q�`�>WKd!*+	�A�q�	�̇uh�Q�+�B�wܨ��xL	>�A�U��[m����s�iD����@�su+��:l�U����#�)̷$��hŎ�-� �m��?b̅wx(��^����ű��Z�����F|�C���c�
zc�� �O?�b_��x?�0�ӌN�$g�D�Α �x(=�^�}����}��\�gs��6�'Ƭ���v��������s�e�?H���3�n�Έ��Ԝɿ��6rp�㏆ޗ^�)#�{U�3�65�(������7<J�'�G��M��w-! �f��z]�~���(�?%>Ԭ�e�0pe��o�w��Lz���t�4��hr_#�ÞDd�w���;Xc��~Ԧ���!vJ$J��x.�:�ڐ�ń��h��YQ��@�,Z9�`�3���]7
a��LCB:���_˭ŔX"�}X�I�lT��&ΨK{�ܒ���6�'�
��偲��f�Z��w�g�d%|�l�U�Oݙ��۷s�ho�-a���w��Tk�1;s6G��.�^�9��n� ����CP`J�,���S�*I����r�rN�P��w��R(���\�%��J�s�.��eql�<��S#i&1��=�KzՂ1Wuq�_DxxM��A�3�ɽq�o���\�=NU�^��[�if�D�uR�\`�6a�\I�gP�A��i��י��d+7/i�5�F��Cd�M�".j�JwD�������&=�%����/qQ�.��jJ���Ղ��X*�_��X�*՜.]	����/�]m�*���)�S���E�������e�9��b�Q�3�?:��������_���F���km{�gr�G(�j������x��4t��`)i�t�P-Q���c�U�떔p����a�q��{VWn���K�Ծ��  �&.c��h'��� �}�%�.��h�Њ�NKv]���5[t�A `JAsN�֮Չ(P��x�G�D®XZ�v$^�r*���Kn7L��Eո��T%J����f{+B� ���;"��y�f��P��+E�޷R`�s��#C)�!m Ov�[;��:�	�p+�x�߷� Y�
w[ӓ�x��F~�mq9�3^��a4��r�L��Q/Fgh_8�@L2�����ع�7;��Lf�Ym,�w���a�fQ#���?��y� �T�Iͷ��]R�`,���=erq� �Z�)
�����Z��Xt!������0��1[}�"	�����&���N�h�X�Ϫ�%��d���Ը��۵�r�߄RL���ue>=�A˞�M!��]*`K0M��<��Q��s.��K��X�JށH���p�m�Io0���i���v�9�ܻ�d3�^S�z���f��W�M�uH��wMW�%q��U��Vq��:bZ0lw�`=[�$1eTf����+���(j5U�iv�'J�h�%��\ ���[{Y$ix|�=����?/�鮯����q��A~�6:iHfb�e
��$��3���u�a�(�:�wv���	瓋�}�ɰ�+j¨�$�NN��w|Ւ��ƨ�r�Yc�,*-��g��7h�+���DdA�[_��H)�L�ш�臰ޒ�	�&�ۂ�s�ξO�9���6�iL%�	���v����js�1�1>��?%�k.�lW4��6��1�*1�83$��Ë-�"�
ߙVC��K�9�-��A����4 �W� =������c{�P���!C2q��8fkn��AF��`0h���$5vu�l�A���YUvȵ��bYC�zB��[���&�SEJ-��m���@�!M���Qs&���wy�3|�$M^屬�=��'����,#<��B%;	sn�!^�TH�\Q�Il���"��C����>"��3��^$M{�O蝿�|�K�ə�dO]���P�1�����n�X�x�_���*�ؾ9J+ю���(#"R*��F0��$��x���Z�ro���|o�u0���=�P?0��^��㣅���b�b^�(�������$�V��Z6�uc`�I�N�,U�M�OW0f��C`(�\�j�(X�3v�<"&�8��[�yS:�j�Lj����p^���%YUUJ��_k�ݲ�ada>˩2:��{�vv&��x �f�*���c���!��������q쁰V�F��O��ґ���Y��3�B6��A�+U�a��C^4�1��:*GG�����=����' �|ǯ�3T�ت��r�d��K6a�
��ӊ 	O�n�E�������4���U=�ȍf��L,��g�+.�_!�Jdβ~��嬆٭)�t#�ˮ3�B��"Ma�LJĵ�AH��=��@���G�(�s�tg���9P.�Y�c�l����_����=�{�UǦ���~��wG5;k�B���@�EH�S����`�P�ԇb�oIv�G�b�G��1��y`�����8�
*+��j�P3i�<$8(�/�a�A���q,��� J�up��ұ�{��6�0#��-�\����3c����2e*��n�L�t9��,������n��eTD�T��e�4�Pr��:��6wy����H}�Pk���+FdѺ���`iِAIem!�L�S��2s�aA�OJ�SZ�٧��[�u���7K����h���8��j$�4l���\u-�Ұa��C�cV���^�L�'�ҽ�N���:d�����V6/�G �4�+�֡�6�h�S�IJ�l1�ͽ>D���yB��|led���	v���ntS ���7�iq�aS_n+.[w�ǻն ��4���E�^;��K	�\���8��Z�cŰ��A��t��4i�0rDe��k JoQ�m�{�x�ˁ�$��k巼��Y��~T[�����E=J�+W�w~������ƹk�`.[y$� 	}E�q�>n_U�iz���T�B��~���8ŕt4�X�u��p�����#R�U5#�H�F��h��#�]��XR�>�0�Fe;�M���9�:wH��b�$��M�A�T���������FX�N�>����v���n�-s6m��xI��@����9��b��[�oƗ�{�H��Y7�.{���HY|{c�x��?J��)dG��6�����x��h.nR@,3ߗb�!���+�|9��S�妨"���^�c��!�b �4M{�^���WkiX�~ /c��D�n;x~�)�R�0<`�$������7� FX�}.��:z�?\�ؼ���k�԰Lg>|��Wt��c��~	H�&	㙗zg�ɉ�'K��É���b6H�L�#]���E&��H%B�&��)	_�D�mȱ����I1�N��UY�->؎������-Kn�m��;��� ��F4���O6f����ИU�r���~�n�xL�70��\�����$|q rKh�kH�G�s�Jj�!�]��tb�s]4�IR�;���r����Q"׎�B4�?}�>��ޛ��G�D��j=�W��v�h�8�
�������sJ$t����U��e���w����w��M�����^�	x3q���Cj��/_�QH�d�I�9�>��[ɼ-�Ϳ'�~,R[�#�h�8�+te��c25�L�&�&�;gH�#G�w�d�1G�#�@խV��c\���J>
!i`<�����<q*��v㱧�f(\^�������}�C���E�⥠�����],�؆5$gW�\D/j 7�8}K����8o���"޲!�9��o�~�Ʉ�����	�0�!��c=q�{3��ӝ�2�n70*��yJ��� �M�h���f���\�M�HV�����}V=��E�a�8�rz�0�hQ�
�������K$ �8����Wa�Q�.�S ��pp�_������d�]LP.3�4sr�EP�2��̭���H�EZȥ�6N(�u�[��2���%��ؖ���##Q{���Q7wsR�G���+�񸀇h�Ԅ�Й�D^܅�!=]�r�<ޘ��s�Q�B��V��Ѷ۱Ӷ ���-K8����SE�a�휹�*B[Z�`���l���06�m������T��$��1��H8_�
뷽�|�:c ���I9*|���9�Ϛ��v��-��B�.���K'��W�~PNҞi�Szj ˦y����a���fYs�5ϯ�*QٜJ�Ϟ/Y���������䔁;(���SS{���4Y������w
µl���L'���v9����?�?L;m��a��A5��� �V�l,�>�|�3*gi����e�"c.�	��R���D��n��.#����LZ&ۨۢ�f��{$�5�a�k KT0��	o�0�U��m1�(�Z&�F�U�(G���!��Y��ټ Q �8�B��DFn��z#f���X6'��2s��e�PZ�[�l�t~���Ek� S��4rZ,"�"���+�u3խ�n�h ��p83.@
�,�n����B�c[جc�=�J0�t���l0q�23V�� �{�n?�4�b���r�d��r�,�����_7�!���#��B��eq��3ӏmz�@��*�g/�Tю]P"`4��b������x��5<ai~k��4Fw�)�Z�x�U�Y�4]��&�.%��c]�,��v-�4ɠ�θ�^k���Z��}@T�����y��iu�K�K�,b�1�3����6�W X��m�a�:Q���N�g
��;�9�^S3_���.s�7�,�6F�4�ϸ�i<Y�5xA���?����m�G�� n�I��(mh�{�����36�9�OZ�0�a�Xz"�<Xw���7��PSFZ�ʈ	s�9p	X������8�����G��VDO�F6<Jx�oXC�=�	�k����jy ��g�H��`$˝ӜƵ��9��#d�J�b�b�a��GQ�H3��#t}ڛ��*�^
�,����ڋ@��n�$2R��xI��Q�#^��u�yIx���n&��Ƿ�?J_|o7�4���o=����ht�x�u�����~3�թ�J����@���e�"Ӡ��E��2�~Qd���Q0��[�F�M��Y�
$���]���?2��� �����j�8�k����V6}�99��qA?B��ڣ��Mn�^��8��ւ �F����"ݪ��|��>Տ~�B��(mc�/19��/`>t��BN`}�QdCF$�8o�yB0�E����RZj.�I�*T��� �X���i�x`E��y��r�rT��)M���p����w'�~����Ճ]�r�b�v��a�\�78w��_�ɐ떚�T �F@E�DI����W�]�[t��h�k��c�}ޡ@U��	p2lU�Ի�DaZ����Eo�{Ap��;Yw!k9C4�.�o��fƴE�, �p\j�e���p;%���ÄߥaR6�����w���YL�xo�-�խ�CIr�ۦ�J�F��&r�O�Szu�S�VY{�P*�R>�ǃ��]�8�b�'!���g��I�TI��c�,b^���'�_�Y�z�Kw���Ro�L�����!�e��Xp�vʹ>�L���]�$�k�`�\�V|%�,���.�Q5?+�a��u܉t��i�Z����t(�U�#_���̳ �b����h�O���b2Q֬��T
u*�3\��14��}��*���J�y�w�[�Z�r�U�|�3\�p\D���΍��o��
����ڰ{!�Ŏ��W���F�yWu%���^�t)���6�wǪ*����UH�:-ޮ��&z��6�&4���݊l�ë3�A8gܓ��M�+��,�x����`��4��q*�U�E.nTe�%������ױ�Y�Yh��r�%��0�(^�!	/�Y�m�R�@�����K@�$��Ø���v���Lw_�?vr�*�v��ݼמ@�����ʹ��<���Pz�ǆ�u�#�2�h��d���'�W��}hݎr�t��Uf�NY�x��p��0���%��:y���
X¿��KF*��]/��,V��~�Q�ل�'@b��NMi�rl����<��3xn��������.����`7!uٛ�c���PPP�-�d�Z-ϕ�%f��זy>�1Sj�(I.^�e�RVXSY6����g�9�l�4���f�A}	��h��d���q��s�ռS���O�ŧ�	�S�On;O��m���W*�`�!
�E���#�&ʚb8��4_m�r���P�䦶��m��E��i��w�I]\1��xu���Q,�\-W֎z\��\��s�h���N��_�=n'�
~��A��S*q��GU�gC9R�IpGP ֲ?P�<;nxH;W���NW�ŗ��[o� �}��I�
��m�����)5j�g��ffM|����gff�������""b��R@�L%�bZh��/���,0��2���^CP�́5,Y��c� ���{.��=
�����I���a�'�	�1%���oC*�d&Z��I�L��*�
60j�Z6������mY�|�f�>�|��N�Bh�>I����}5;25��	/��X.si�}i�h4��A�7�!6���>��>�!��>��=F�2��7Bx��l@0�?A���>�2�i�̤�z�"���+5�O>�8��i���V�eB�b	�$��ꡉ��?�'��̈T�ܻ0��<�6AFwDY��T���W~\�/�1���T��qp=9R��0���4��#���o�ڻ��2G^t=��V�蚣S� �r��_l	�,o�� ���o���x�ӎ_�����Z�n.2�j���Gp���ۄ�"�T;yޛ�G*�%��Vq���p�\"C3Z��K�����Țm�2�	2o'�P3���6(�A���j)gN�#JB�(����7�5�Ӑy�U&�!�_���R�=oNqZ��P������Uz��B�B�����ՉuR\�y�|  Xe�O1Hj��Bh��Tt-���%��ީ��`�ua?�h�I��3�u}��I��k/��V���X^�����x����.<���yЏ���qn���@m��A�Ǻ��E�� \î�䠸G���k.M��&]�)��f%����$=Gl��.�33�ݰ���Ҡ�F�8uz�W#)�7� ��k<����eh���1�NBPr���Ƌ���ĵrק��zcM��� �Ńj#	���r��z�Y�)��ܣ�fջ�hU@��b[��#�xY�ewf�/�M�Dm�s��x�ښ�1f�җc�B��g,dɉ����F��A�&���a���C�?�{ܠ��\�F��P)�"��kx��Z���i�77�4T��Q(.F��a߅����@�ӛD�A�����,O+�I��Ö'�0}'HT�(*D���L��������3�騋���-!.���z3���}@א;��zB&�p� 3�X&4�=�]T]7.��馅\�XCX�2(VQ
�[e�	��}�N�&���E�{ ݾJ"E�e� x�����h9(���N�#��<�1?;*,Ͳ��īli���螢�-���J�_�ほs�����䐇F����`�Y˪��;��OC"	q�w 7c�;9���R
�$9���?���X�q�3R'C���z��s�v���	-�$b?�O�*����D�q�3��f{������%'l|�kU7������¡����ݔp<+��4ٽM�� �W��^A�Ǔұ4�[�9f�R�rQފ*���<Dm���
�M�5u���ܫ�"��"܆vo��hJ�DR�ߨ �M9�:݅tMBa�T`Gs*{m��)�di\�B�E�Ӵ����\l\,�C�Q��嗼k<0�C�[������ZE3K �݂�;��E]�"�a�A�^ d�l6�� S�CRp')�	K����X�4FH	A���$������Z-v���/c\�|�d�1�O���|G�\��<�|�)�H�ӊ�k\��l��z�!�Pyt7��{|�pG�/��O�
�l��8���Alb�k���Q�\X1ḩ�����`���0��?�ܫ���(#9�N��77��@(���{��a��o]��U��,�Eg1�וpRdF2m�"�!���)a���&8�- G�-��D=
U�et b�0)���rp�|pg�\_��s8��
�g�A�g���Q�2n���ws��\���J�r����\	9x���4���.N��*����������:~`��^����J��<5~�X%[��
~bI$��9��޸��x2�%�w�P�m)8�����%w|��1�/�c�VH?�<�r&΂����*�P�s�'�!������/� ���r˯�@�{p�S�`��܄�+���b�J�m[y�kW"v�����!��V� �𦂂�)�43�L�]����=�x�,��ʆ� ��_�d�4����ô��#
��H�r*��n�+�f�^�^�Te@��I췐L#�0���I��w�b,m<�8�Üj���p�=��2�s�Ap�(���u��棚�����lE��M�9*D/��VW��"����xa���b��	����q��Q�J�rю��|�B��
j����8��.���2t�O�ku�@b�6��%��?�Ｔyo�ϛ��=|OV�������F�"����1c9c��4=��k�&ۚ0;0�)��,,~��;�w5�;����^�ek��zl,��$�M]P��8ԉH���3�o�Tʓ�Љ��+y�qyxL���ٞ�Ak��O�n�C�(1	�.;޹q|RyU�;i#[r�q|TwJ�T���:��?GՁ�>V��~����.��_���c�W�jO`C �D�I.������� H�[��p2�E��V��)Tʗ���h�LR�����V@;!�?�:<4�j#�U����d��X�I�0b:�� X*�gv�����B����j��N4�dF��@E:��e��ҁo**qUS�z<�!�98��u���D�J��ܮ��V�zڟE˥���>షs�1L�`5��V�	>�Z6G������bz9@�Q�ַ�֧�}u��i$ ��OH8{�n<?=�+�H�|�s�ʠs`5}$��0�}��Wg��X�r`��gc$aDO��fZ�?�(ˣV����-���j�'%��2~�"��\�&���t͠x&�+���#=z6���ux�}r�l�,���C��!���S.3<�m�!��[@�Z=@�}�ܬiR�Ѕ�Bq�'d���T�X����cd�lͬ��;�!y$��U1�+kE��_���!�����=��N�ץ�Z�p0��(|�+McA���A��2@@�V���YT����R�^���wpȎl�mtMm �vP9Q��>�����fh������X<̎��B(����L����*ꫨ�(ػ�8� K�F4Q��������3�# �F����F���PW }�G�G�y�,�	d�:PC�Li$뤾�-
P�T���_���s(D�VmR{?٩�n��g���i���S�����~&�`�-�'�0�M֪?��=��01��O���"��V\�����z_�7���i:����0���^$�@s�z ��0�A�]r��MC�����6BQ�d2��|��u��o����3��a2��Y��W>��SL�����m?i+*�D�uw;ηd���rR&��p@\k���*aQ�e<Ȋ�}'�\�pE��$0l���c\J��[��D9�,J� O!�18`�A��g�ە�A�|� �����]_~igA�3�y�،US��C���.l#�mr�%G��s�Ql}�2h=�-�z�'�y���޿���}�?�b1#�R띸V1�)�u*����묰e��۵,Jd�3x�J%UW����¯x^g��~H� �B^�u�_Z*�ޅ_V�9��dGp?���i:|�&Ⓙ)�Jw�J
�� �{�f�.���$�6ˋ]o_�]�e�)ގ�#W��8۞��:�L�IӾ��u^<����޿F�H�iDm�9�k$�Z���|���T��%H}@'$~�_��|os�[}7Է��t]�����=�i��y~� :�������I��#z�Oޭ���\���v)ZMqA�����ȉM����Wg�͂��3d�d%�4X�� �j��jMa��ؘ�d2�U�/�qn�5��/wm<c*
&���3���@��l�.�q���U����[�L���E�C��_^%��0��y(+��*7��J�i6tY��C���B�3�fSͼ�����=b����gX�ɉi�G�q_;���:�l�I!6ђ0F�A�YK0����t�z��t�K��Z{,�C�c�.���������PX�!��#�[��1�lFJm���m�kS
��/K��]jR/�4���-�N�Q��>�e1fk~;���S��+N+(k�=����}\�HU���q�cb@���5�_|X���r��]R?C�W�g7���r$�<�%h�����cG>�6,���Lc��
d� ����i���R�`���)cӣ��\i0�̨�� �6J8O��R<�$�&��ĀE��m��L���k��z���1��J���¤��ȸ�������i��6WTg��n$�,��(�߇���;��ҔƲMa,����=��f�jK@שd3zw���e]��j�d!znC_�\���܂������J�lt�`;�Z�h�"��Kn���礴>��4a���\�&�!��)��x$�nO��$tx��tO�*�ܯ��J ̜!q/dQ� �C�'/�W�)����T��fW�� ��!*���lE��z�]5h3���||u��5��<Yo�I�����Pi�k�-��;�t���5y�A�����.yD�u�0�/����(�������M�^��`8 ]E(o���%p^�b�.�#.9h��OU�����O�u�+I�=�<�t9�㇙sa��ΟG��W~��X��H#�HHZ�>�c�8��'2���d=j�Jk��dlݱFViu�`�y 1 �Ԋ����)yv
?Y���(��Plm��n���:�-eP6�2��@fC)�K�����YH��yw��{'� ��1�4V��7���Xa#�>���QdnO�Ck��2�gWD�	�w�?w3�1󅏕��AR��$D�K_¾Ȝ��]Ο/��Gm73��ԗ�V��ZE=p��7B�i/�wa�%�!�zU��k
ZƩ������Ec�O�26`��'j�"G�w�7핥��뎠�Lfg��@�����Uo&d�s	8���?���;����t{$,�t-��'	v�DaF�x��}��]X3���$��S���+6}�_N��u�7����o��i7�TV������;	��\׋,��Ϗ@���WU4 ��wUn �2�6�)�4O�1�=��C�TF0yV���Ԏ'�����C�2�,m��>^lR| n�m����a��+tu�q�0�l��F� �	Ev� f� �J݈u�9�$��*_Zwc���N���:�"���mw1ÿ8���n�V�j���
�P�2��"B�M���gk�����qh���[&��%*�����m���R�Ⱥm��P�d��@�����O�V�����)*ק �1r2�Cg)�h^5����9�2�%�k��_���F�����b��+i��3�㢢����l��i��!����ZB$���΀��Gk"�k�.�^���g�}
Xc�X~T)	�^_�D�`��/R��ʻg()[��J>�5~Oѹ��Ĳ�<<v�=[��`p�6���Q�M7 �n�_s��ȇ�)��j)��	�M�y�
�|�w/�����*9�ܕ�QY����t?䚯�:�6��G��OF��s�����'t�P�]����	oY��6A�E}z$D�X�^5��;NF�N� j.���ț��߼"-l�`�Q܈�� �%̘��hj[d��!�9'Y������}Y@�=յnd9[2~�{���*ƀ�뀊�=�X�k.?��	��h@�y���
�:�L�F9w-^IFu
���Zy`Ƚ�z�"X$/Gn��g���_������8�$�c��l��&��!gb%���W�kc2�g�q&dd�����-K��l��W���	�D*M�D�W�e4������{�n��5��H�ba�/˦/�/��%I�������ּtL?�
C�~�\r���O�e��5����Y��j�����JuO^2�1�~,��׉�L.�Kcu��`��`՗�@z�:E��O�iV��lV,�Wt;�L�j9��AZ��4�vɻS�02��m�Ճ	j]�B���r%C�?��V)���8X��^`�R����Ǌ�4���b��>�k��|�����9J4&��COSq���k@n��)��	<ك�5�ҹ�fwLPF�j~eU��T�lO	+�~�~Qu���[/�E�w�UJ�oyyJ����ؒ�sA辍�k������B-�mB�
�5�0�	EV!:��o����c�����P��u�~��W��G^����x�OϹ|�C���a�ucrܺ��G�ؗ��B�#1��tƑ�Z���jAt�7�i�8��@Ol��;xD��xHX;)���� U�C�/b mv���s�.��{)��C�_�,�SA�7/��������W�K�Z׾� @X��tO.Au �`��� �bG��Gm�w���q t(�_�]�?��vx	r���M���.��h-sZc��Qz��ONK�5&�g?DdFu1wK�ߒ��q��,�����oe���]�8�9;\8p�E�{	�U���ȶ1Q
j������t`�ed�l>iT�JS����\2������}�J���
�l ��w(WC4쒭�Ň��s�g/+���1{��y�r�%���Q��?�lFR�ҟ��J�#�k�q
RqaH!b�����E1����e͝�� #��L��!-ac#J2n�oysyr_�eA��`�CU��ں@�{l�Zj�L*&FK���%��""����ǟ���� ���+~�,�¾-�n��~��&mF��\)���Dq�4��:(�S~�P`oF������tƈJ��3A�����(��F�H ��1����UJ��߼B�7��bU�ַ��ga���7���`QՄ3�6��Θ�j뱓�*������snӔ(�ӳ
y�j�#�L���|���̊2�Em)��W� ����Y��7��z(�Y_�۾a~ۂn;�W�Myؼ��8u��2�l��Z�|aPU(F=��ڕW��N���	�D� v�-)`�;ѢPȓ�b�ڍ��\�U4�G���C��f��dt�8����a���.�)���Aؓ���#�GS������BEM�:��[l�#�ANr��g���.�C�2��9!
����(6�ǝ-��S�[�Xt���k��AzD�q8��}^a�����#qt㯛+$3��xG����S�kpy�)aP@�So��nG��k�gu�s[֣�qAw��� #=WT��3��/B��3�ʁ+�Ml�m��cp�EO�0�lnY�K]]�b�2w��ґ���?�h��8Pfaspt��*DR ;�nGs�k���H� L�J��ߢ$���'��@��[m�t<�0�Q�馱�E:tes̈�B\���Еꡅ��i���ū_fsӈ�Z4&��v�����5�Y6`������;� �/���G��s̈���C��(��\�n�u]9j������3��ΞErMI˓��+�quM���=WS�4ߊa�e�z����cu�-�k��<C��ʫK���/v0`�Ӎ� �ݝ��z��f��㻇�q�ߕȖa@Έ���arkĔ2�L�O���zYxe���X�N;|Qb�4������b����o���q�hvtJ��,XI���B�T1�ߚt 
b���nm=r��[�#C[�ïrR��)$$Q�Sp��?�o:i쒵������RUn��P����w/6,� A���h󬆘�Q���L�8���\��\���x�1�~"&�tы_,O��aܠf����U��tps����]�!�N��M����f^.�f��^`��XR����I�η�".]������+m�!b��ߜ�a��_v�a��7��1�`W�I��=�-�֓眑�@:yU�FQ{T�dX�E���Z�=�m-��Q�u�X�L���,��i����=�^b�M�iW�fR�y؂�n�u7e��_�˷Y����4�W6�������'f��R�m��P2�w\�l��$�(������^
4�	�GHi�T��U!k�<ԑ�{� �יsf?��Şm�'C0�;�m�������z�ͺk���Y�9خ7l6��;k��a(������!��CE��w��ح^�=��ۙ��� Z�����P�׈�~�5��X�t#��"�W�0�mHJY�z���F6�c���
o��j�IR�Ǳ�/Dݜ��zA�
�����4��G?�`߬V��RtXD��Bl~�n(:lt��W��O��aާ�g���%��H���,�~�+[�Td\�ّԀ��̃D�A�Wgl��:��M8��8����ȝ�]�s�+;f����^�B������_�\:2�I�'�0SP��eYp����vwG��ah�~B�4l��ʮT�t��K�_w��#O���{Vv�/�b��驚���l�=Q~H8u����xs5'Pi������TN��#�~��m	�#�q�玡���7�;�R�#p?d8R���I�ԍq��և�uz�萊�d\y��H^T�wF܁v-�&�\d��=��9_`ǆ�Y�3���|{�c.�8�6;Qo�����[����v���F���f�j��+k��8�X���C��c*5.�55��Z%��80���S���!B{�"���$�X"�T��w���~<`>�wyyd��,f�I���h���9m��UM���n�M	��^��
pW�M�G�{Jk-/SC
*R���|>�~[�szwj����A)�>��e]w�+�V�ԁ"^V���H�K�������X:�RH���#��3�$�?��Q�R��u��F�+|�E�D�*�m?2qEi�$��gf�Iu��껭�"H���ӌ6E|�;�����+�>uy�h���u�7�ʙ��3ʗw�ʓ�}���F��I�zC�o����'�6��/��1���+�fD{4�k���=��m�ʍ���I�=F�'�:��e��q�V.ov�O���(�h�3Y����c8IR��5�+�`4��|��g#��ӻK�jm�4��q��6���!b� 6G����	��!�1�C�ĕ������i`�U*�n=T}�NT�·��P���$J�Erk2�cyJ����i�'�x�mp�;⨓x��m�<����u�����Eä�;� [�D��N�H)���&!�"�@h��]�u�Zdgߥ��/6�qwKP)�K��NL�5LcDo��MhBM�X?����bH0��u���-�x�㇈�]��KR�O�>;��������c�����^ՙ���y� �T��S���+k���R4cc.�P�lD�|�t��9�,�L/�z�6H����:\{7Xw�k��l�D�+�/�e{HAF��0=g�gO�]"��|``9u�A���]W��,��F�M�ٿ,�^K�]�ȗo��n��c@�J
�P��C���b���%��6}c�kQ�%�p0��rA�3!}�k�!S;��&��@��.6Y���m��M������� pvF�����'�.9L	Hkю	S�������k�z��î�Ҿ�k���c#T ���g���|>� �ؗAN��l'�d�;�@
��<��|�i�&�^����1\�)��y,��iqt�jA������
X�oPC+�������f�0,�L�ZL�$g� p'\a���, ��\�.�R,��<��q�	^�F�Q�4�Y�>�{����;��C���~n΃>�HgX;T!C*ס�ѫP��-���~W�V6'�2���i�-��$�T�.��2�E���;-���a3(���5����F���k��u�T�@��_,�&��]��W�_/��1�{f�wW�1T��9��F����'�bql��$)����)�S�l}��8����ěо�(�A��A\P���L��Z��|��H�\YO�sU�u
N	�_�΂�T1fZ��˹�Af�x�"9�>%�mq�������S��C�̓��)l��p��lI�+$j�|]�98�3�L�ox3-��1C`�M��/�y4q�)�`P"�K>��S%����(���=�Se/{�sL�ڗ76��&|i��ᎊ�Ǳ��|��/�wWe�$�~�(�V�àh�軧b4rym*{z�c�� ��x�v%-��2}Ά�w�I����PL��p7'�7v̩Q�K{�'�\pHYW��S�BM��LC�?��Uz�G{�wR����/�W��QZ0��� �,/p�΀ ��g�[�V?{�|F��k�ij�Y8���r/�~�t25�xv��F̐��g�{m��ѐ��o'�b�E�/)_��2M�n"{U����v�6�l���F1êl�+����b%�>tG��H��e�"�2��RD�u���kh��H�}t&�K�X,���"%�w	M`��;&�M�����a��ԅ��!�/�d"{<��n�ګ�M�	�rt�pY�KUHj��^U��;y���p�iRo�VTmd��Y�g[�m(2z�a2G���C	��y-r�\[�PMV q��h�`k��n��)ŊH�� ���y�9�<�H��$�*�*]$h�c*D��[����<�|S�N>�y7�vX�<ߓ�6,T� Ԍ��K�S;Kߊ(�=L(%��9/×(v��5ƒekޚ�"n�0���c�+�?5F�C;,��?����(�kd��&;5�i*�T�������x��U(�+E1����0�"�i;P0��7��������]�MФ��ݒ�x�eA�	f�|3	��m�pX����U���dxH:����_���=d�!�S\>5�/6I&m�"#���Aɬ,<:�l�l�j��	��2�g��A��X��'��e�n�p��R�#���G����N(�hf�r/Ŵ��޲e�j�B��
7�����uiN��ջ�!���]��B��sap�p��U���G�Ψ1F�H�� k%���A=Ũ��;�W��q䢳vx�z8��yD��5-��ՙ�fu�[��쿦�R���%3�Ŀ͏O�ղ���a�b9�+O�^O�GAA���e�W�k�YH��)�|�ޣ��\�����0 �f���
br.XU�r�X��9���I��w�%�oy��f��.hAu�xĴWI�d��:@X/���Jh��W
���"��U9��dBz�_��T�����AΘ������o��XF� 3j��mZ�<��|����nJ��ȝ
�6xo%X+�U�#��sU|<I`h�h6%qLLF�;H!�g%�`!Ώ�V߂��)}!b�ڎ�����Úv��K2z�o�q�d��G����1p�!H�vQ:KgR�/a}�D���{Cxb��y ��@W��y�����Ot뇿7�//+^�K�j���*7J�f2z���jʑ$���w��2D�L������7����çB�nL�`��H�J	JV��O�n�6p�f
~:��c�'�Ðu�ԇ��svέ �t��W^��~�
mQ�)��c�zJZ��X&,Ga�M�s��ݝ,CI�yR}o�?�.� �e*:�$�M�.�x^M�,���ӹ3�sc�V;�n'E٠<���3� <'��FU��Shd���*�yȣ����X�3H��)�ߧ@^!k-��j����Q"��"h�*�@m�*�\]Le�X�vA+���餖{p,���ZIUQ�� `f���2s��m���&ja���9g�^w6�㌳ӽ�����+n�Mzd�c�ȱɺ�pn�b��U�3Ԥ�xoi���e-.N���� ��"���@[�wgy�"E�!F �0����d|�b�)���ɡ����8����x����ߚ�^/�N�`QB	KΝ��z����������>4j��c������Z�����~�*Ըt�����ew�k�b���zj��w �r:pU�W�����Ar̸����0W`x�򝛰��tv[M7C%����r�$�_��[�ݧ͵�׏��1�A�R����.l��	p5����ո���>i��d��H���{]���9��o������G�)x�VE~Y�Z3�F�i�����A���s��!�+��'c�jkim&܄�����߷2��;:� M������k���4�	�X���1_��Egrp�J���(��Pt\o�n%DmZ�����W��Ӑ{�+�x�p�o�09ۿ0�.��f��L���(a���wJ��17��ϳ���_�<����:s�ѥ�qm�G���w�`�.Z�_G%�h��O$�iH��!w�hsmlrQ���a�h�����$�Q�z�惴�L��y��#o>(
��VN�)	�������2+���t�/�7F��E(�w��#\YMῳc�RQ����	w�fx���8S��m�x[�l)�cgן��$c�g��s^E�7��tf'R.�b��A���JN�Z��,�Φ������F�+-�4hH$v�3&�x��`�Q	a���{�����6�y�<�rEn�1a��cp��c����c̽긽�X�=�6W���u����`��NU�XW�Æ���9��!ͬ�,���Nj��X���X7SgY
sR��aؘc�t�C��� ���9
G k0��"�t�b(�5���%p�` �P|�qA�X����i�t�x,�5� �}����O�h�; ��ƙޘ�Mw����"���x��z�7N֑c�+�G,�<('q�~���_n�����)�WgLT~g�0a`�С��8���o���C��	�7��.W�p����p]"���W��&�r��8�'v9u����ܜ�9�"�ԱZ��$����D�
!�I#�7�B�[�R���O�b�+
h��W1�=p�T���PomL�";[�3�6 �+�m��f��lT|}'!��9�d��=�X*&��>���2�'���_[�_�q
��He���cϛ ��xg�r��'�mgF1��eC��7�꾗����T�ThU�w�\�;ͨJ�mu�v	WF�&SY奘;H�\�s����bM�_�nT��.�X䄉��e�p�-��o�&�����R���(@O��{1:�F:n��"�"��-��pu�k|,޴ڪ��.�^e��{9��E��0�,���M�Il80~���j��DDQ�m��ec�y
Bwic0�󹌹S�G4�;m��p:��\Ȧ#bQ��z�{_l"8��M�s�����Cy�������J��Ϸ��i���H�W���`�5'Q7
�b�@�YH	��L!�'����ΎB�ۢ�v�L�����f^�޺DV��ߧ��b|)�ܭzl%Ųۤ7L�в��p�8nA@�7�j|�u�
QNэ͜%0.$�I�,�]�|'Ey��Ь-G����;�5+�Ν�]p$f-�� �.��B`p�@k���0HT@��o�* +\xև��tĶ@,,�m��BE7zC�?��2�,�F����Lq|~J3o�0��K
Ĭ
\�G��p�����!�,nX6�^�-.R�@�\� _�C��:�3="�Rp�#p4��63eim�r~V	��f8tڐ�����x?1!�������XSe��4��7�?"�I�J��_Eè����/v��ekC[`2=�R-j��7�ɐ�۩Fٟ_
nz��}7����L&Q㑇�6� ��r�\���RfoG �z�nwJ�i��i�i�l!5����F8�{g|�s6\�w%��b�is���\!���p����4YJ�����m6��dM*���i�a�8�2���9àY��=i)(l�=��zV�aҲV���O�C!�D���X��0cx�	�LQv�g�W]}
ҊH+�O�t��HЊ�%���]���GzD�RP��1��A����#���.q�u47A��4�Py���<�{"�ϓ��f{M�4=�
�qG�������#�$��l��W������@<\����3R2�v[Q%�d���Ex'7��ݱ������ɪ]J����K����`%���2guڗ�6Z������ɴO���Y[��	��F�.l�P�}$�gZ�O���?��F'���&E& u:b@IVL}zZ}�μ�NU����.�k�<���ۛ`�֦�l�r��?y�z�9�p�G�/�״�>�V��ۜ�R�tp�w�,�f�|��,���}��a�w:�E$��-ˉŉokX���7�ͼ>C��̮Hx˶ h�'����+XJ�b;�Yj�������u�r�,+�YS)��ӔF����W2t>��wc::���_�n����Jpo�5�X�{ .u��}��L�B�5�E� ��B��r�@��/Bt>��<Q�πE�����=	�d�z�#J��]�Q�]Rf_Bl��>8^!�К�a�`���K����}w 5��*������lnLF�-�0�viF.���0XZ0V�dd��(��5e(���v�>T�ͦ§���yԌ�ե�v���֛_B��F����=������B#�K޿����_Q1���w�JlTX�A�a��W��7����Tt��e��)��W&�{"߆]�S��1dc��}�,~eg��SM6�/�1�����w��B�^Ȫ�38��8���#��{,i%��/͞��H_������ ����ل4iH�ny[Q��~C���f���QGBb��<%�~�у���6�9�_h�_�o'1��%9���h؛Ŵ�i�����E�z:�:��B�k�\���R�86�g���9���;�����^a�b����u{�	$��t��]b@տ	�����cc��h; �qO_��L֣�M������.�g����������2N��=�e8��z!2kϾ��� ���\�Y��QV�B�8(쿴m�i�?��8��|��������p���	Z��eKǛ-Id���6@�}C}��B��H�u��P�ZY���lE���!GU7J�A;u�
��6�{�=<6sr�=%B������U7|�w�����?�*)*��&Z�|J�ui��i��!.!��܌G#$���D���|wkٞ;� ��7�����4 ����]c��V��a�M�u�F~A�pȑ�SJw�W ������C�9���2�C̅�M���Ho�J�AQ�lM�b�0b��p�\�L� �+Oe�)Q*��y�]K.�PVe�}(v'Z�nӝϑ]�N�JL0���Z�D��ſ�;b�K�G����p@p¶d_ S�m�J<�E�tKZ=�b5WӉP�w��u!�D�G�9�x�e�o
�)���;�Tg q�UL]R-J��U(��3�5CH�W��-'�:**�ر��zl���c�Xd��X�г��]���/�c)c3����������|ǐ����ي��E.�󾄿(� p^M�O==�s1�i�ة�xJ�o�}H4$Z]z�S�'���F��1Wh�v��5kD��"8���,#��]����{L����2�J8�v���h���t�M
8%F�=i��u��������/�Y~��v��Sr��h�&�$��uF���L�Q@��ZO��yO\=%ϑ�;��>؃2�n�	�,��G��,/:��3��:E㕅N�e���L��V-`��4%�'D�y��ij!Ê���f"S1�$َ�ٮv�w\����Oh�������L���� h�-l�W����%��|�:����!�s:��Z�HSD�V��D�=���V�x�퇟O,.Y����M63��Ho"׃둌ũ@X`~գ�f)6�[[�z��?��t��9P�\"�L&���:p��ف�νx���ڐ���R�F��yl��<_e��O�����|~QC䠴U�v�aЛ��yO�ۯ`@<�#	�Nۛ@�d�Sh�oKHFa�
n�ѥ6#�(�c�q��l���S�}�z$-�N啈�����������>|�)�	�}�����]�P�^�xH���}�r2à>P='��ӄ�z�p]-$B�8��M�1i�C�lˈ`�#F�!�F�����D˝'��߹��P��%�"dw��_{6hO���G��j��9��bC|N�A��b�I)Z/j8�t�;���j�bF�B��`�wŧX�t�i�HaJ�n��z����8�}�_�P�����@9�h(�����Mb�Z�p��}�o�V���i�T��*�9AI��@���i���<�L������j�:p�N�h~�|㗍�(¤�=���d*�;�}&\�h=GIw��s��Z����dX:-��'�]4��R��IZ�Q�S>Q�Me�l�(is������Q�l[�l��QF���箞��b=�?�%"�����ڱ����QrA�qN�ʹ��S����D�b��*�]��Km �����h�xM.�54S7��<�Ǒ��QHV+z�X6����݉�~ߴ!2"�r�B�ˍ�I�u��tDK�M��X��d�o��˝� �J�[����
;����b�e��X��M,��$o�4J�K���H!P�W6�i���c��z�B�����2�5��{�)�� }��ޯ��qc8���Y�����u�u|��HA��z�$lv�1ΠIk,@�@��|LaJ���b����8.I�8V5���8����T�X����T���h�U����H>�tPl�;Om�}1�� >�|N�b_m����������(�A�FT���X����_�tK� ��#Z9 �y�����\���rrZ|y��G���/n���WP�s7F��J�ɉ�f)6A��&��/m���l)�U yj+��� H��z�������e�j��\(� P��m�����I:�0<>
�|��%t��t,���k&�"�L]��x�Ts�rƇ2�@q R\��H)���#�"|�o�e�1��Fww�f���Ԥ�jh�G�.�/HH��*6ڡ����v9�*މ	�6�E��{���X弸3�]~�,;6�=Z��o�#�S	}r��_��[J2q]���N��o�lѧL!�V���R�K(��{��u]G���;�00̩�'QA�=��~�H�e6M%nlaF�l�2gp��Ep�
�8;5�Ek��^ఘ��4N���m�p'�R��_�k�4�E@��`�lU�Zxƍ:R�|�z\�;���(��L�#|繦#9IF�Fx�+��PǢ�{�oo�ZB*��&���s�@JH�u�2�;�Q�W�j�d����X�X��lkx��H��e+���䇸�Mͷ�.�WhF�Nr�G���
�8������w�@�A��tȋ����gUٞ�))*IDGwS��҅�y�ͺ��+�P�V^����E"���0:���B����gD�L�� �ǡg����f@q]�^���B�~yat5�x�X�P���)�J� ����Q�B�;o�7������9\e�����S�������E����O�o��c�6��/��1=�~��-n<�b�©i��3r5Q4)`#�]���O>����iRL^������I��J��i��e�@�S�����,�f�^VFNh֖����#���NA/����� ��5��n<�l�ܽj��!A^���8��H��hg�9c���I��q�Qa�(�d��N���=������򗇹�8�3�l��)��ťh�0��%�#��,�g?��ٹ1���dF1�|����3��b{KKHr�`~-�$�� 9��s�ï���c�5�K(�LcB	`T͍pB���[/�~��uB)����O�rp�S�G�dnaK[3�H%����L:�~A��*3�_o _��Qd��Vg�*s��	ð��5���>)����3_��P?b����D��i�u���"o��yN����6E:�C��ڄ��պ[Ι m���A5/fd��7ݍ�Ol�����Й�7�`	��H�+\�����f�sw�q?��H�"+������h�1��Gz���G'�L�L��O����s\���Dӳ��ݞ	� �7PrY?mt��Yc�n���]����i���9ɷqY��>��$��md���|����L���l�tT��+��=�<�@c
�v:K)�k�<��例jj(�$������Y��q	<�V��{�jc�).��9	x�cG7����CI#�kd��pFX��=�ױę/D��h�#���qy�8n��I���x&�9���X���u;�w������vڶ�t}���U�D��P��9�R�!����T:�7}����䢿��}�w�����Gy�$�U����7cޝ�?K\BGPE���}��`eJP���]��2{G�:j�V��h��dZ�mO��>�eq����T4&�+��µ�����h��M�[���Qb�T_��J�z�����25�fi�YG��R�?Z�v+,!-�afh Sj��\T4)�;�l*�.��q
��i�0�̓5{y궅Ը�:�.̕#�I@gG�i"AN;7A%U� ��s>�K�ǫ"�ň�ο)1,c�� X')֠����'�r�C����������K��J�#�9���U���sK�?�U=��L�Uz��c�������oI..a"Du������s?va^����Ɯ�䏵<hC�|���H��X,�$U���H���W�G�n2�	\�du^;P���Rb�)��y(�X�<ຈ��~�	%S��u���/,���>���ʙ��5+4]�`�mH��;��Sw+����2���Q�f,A���捾����=3��|�8z�5�i<��_�}=�S���ѯ�}W�2W0�@�u�h�=���K��_}�b[pO���	ܫ�YS8�p�<��8�?+��R���E+o5��C�(�����5E�.�BI���ZG��pҲ�>��;�s�k��u���]�8v�)���w��MY��w@ns��?���4�AT^$>M�Tz/�V�uǪ�����C����[,��5nntt�g�Z���G��{����c���z�}�O@r�� XӽC�{�9��)� �ae@�	(���%p�����j'�E�3fb���xW^��d��\�GBs��r}q#������:��`c�]�a���w������7��	� ��A��QF��`=�z��lO��'b��u�9�-��R�b�T�+�,�@��>�l����`�
.�H�3螷.�xG�ߟ��U���nҐY&X�;���c٨���j5s`��KS��b�tP3�0�:����yļ���l�a��:lӲj?�o�X1�@t�)5<���jl�C�8v_^.�<�L�(~h�����4r_8ʍ�8L쀃K���,%������*��v=9c+g�U	��Пj���T��p�m�/_�p�%v���s��^�zU�&n�f��t�]��⫡��hcO?N;����|�H6�(zKR����`�7%l��G��,�(&
M�A'��O��Q@�{{A{�����ݡ$S>���H��D�М����w�-}m4�U*q���� �r�X[NN���������玁����Nh�56L��Ծ|��R�08��^h�Qp�KD����[�{b!��}i	�O8��>`�O*w�A�Fm6O3�؏Ɠ~{9�����V�Q���X���L�ϣ�ZA���2�6�BYZ�-
�=dE	h�8�qu�5|�wl�m�j��+mu���J�\�+�@��K�f�0�C���{���aP��n�~'>���t�ĺc�T᧊bז��[\D��:S�v�.�i.&2�^�`�s*�֞�} ��&�#R+��*���D	ǤVK���K�6r��-9�['�+��z����_���,�Ǿi�M�`G��u̀V�][�����Q5�)OL�%�Is~Hv���m���"�|?/#���[M���r��(4]H�Ü��V�
��<���6�˹X����~����N�҉*;wސR��-��C��&���b�@�⽄|x��u�+�bA#4;$>�Bq=�0�[���JD̋�l�kW��bV�zb��hUB��#�G׀���S�/+3��{�s"�xж�{�@���EM�i���)̓�R�T?�h)�� ������+[���FG���N��&?����u>=U�����*t>�R��a@����� �.�d�. -E߹����s���P��ƥ���be���(��x���ʖ|�.��6fh���*�,��`�"�5�S�XqX�P��3t	��a�7�-l���䅻���)e<�}�qЄd���D ���@M���d5%1<��m35!Y?�۩�R;�غ)���}ӈ^�|�y"h��6��Z�v�Hٯ��6s2M޴����Z�ִ�c���R����n��ך̆e��\j?��0��84� �� ?�4����M���G�} �%�=T�;�F)��Wv�RF�c�S?S)F��%���Ā&wj�g|'>�^,�buF�1A�qmY�����E�@��ysM�Uڝ�D�Sd�"����2g�Pe
@�*���70n���CCD�옦c���v#4�bk��0��W��-fĮ��.��9���_���aw|B����L�"�m����������7�|��5��u!9%�)G�u�����Gcm�%�Nu*V����|n��?*��'?����@���x����ˣ�N���\X&�&���Js���Xsu%��Vt�,;%BF��)Кmm�f\��?K
����I�&Dݧ���Q�ЮU�0��?a���lv���(w|F�5 jܗ�����@�����v!F�.�o�:*E�+R�⽩�Q�� cW�#�V����o���:MQѐ�dtm4ޢ�w��)}+��|�oR]�3J��k>[: b|�t�1��E_�=�$�"��� ������}q��@�1y���+����]7����,:�r�w�,�U�"�����8+k"G4P7|$lC�4��"�����,(r�@gQ���c0���mX6I1.�j]��`ĺ��@�b���''�[���2����t.Ŝ�T�� ��W\����dx�Ňʩ�S*K.�	�ب��M�iKG%�<.�=H�F��ֱ	����c�m����T���-M��±�,K#I=�뒐���bNᙊ��ͅ��o���C,�=m��tZ��hK��)�'^����̧��8 ϓ/W\�aL��Ku�����k���F8\R����x�m�ψ�CC��w-8����k��E�7PL��̬��Ƙ�9���[��%�~r"�u1%��*��]ť�����(�+��C�33r��==�f��p�$�wtS��{҅|��f��G_Y���0b��"����S��&;#b�.-��d�cOy��uD� }ɣF6L�l`���Ď���nQq[�� tC�ݬ��$C���U�W6�3�)�HuͶU�#��]�x�{ϭ#��[ӵj��t_#�/8���i�/UB�Wl�1�&���y5E���$�'y��3ga�2̎Є�T�_+5l�Q�:/�W?�	������ǭ�At�"���ƀu�g!�F��N���ov���X��ZN#��[x�}��)g�v?�n*QAG�'�|��F�JZI�Ȑ��k �N�R�/�9'��;���z<{��� ���x����#}��=�D����(��M`�t�.�Y�u��k��ǰ0���3��o���3��%���2���[|�vT�-�>�"��*���"�o5sD1���D'�2~k���ώƦ2���I&b��7��J�7���^�J��;i�^��7Y,j~��3w��.�����~3�]�|��jM���j׭fi�9v��c�S�����ǆ���MC��C����
,@I�V�Rs�����T���d�d`�`a��H��`�4���&��"�ѧH�T�G�����68���zR 1*�z�����c�����|���'��\r;E�R#�ř�lTEs��ӱ�WDL*����yŗS�k`/`Z�_&w�zҞ`D����f&�}�"ϟ�����QY��M+��{�C�e�o0Ż��¯z����~^��A�Þ3j�zN=��U}�Ge�4����v�x��H[?]���V�l��"�P���>�w�����)P]mѐ���H4��8r�`}�mD3O�W͡�6���J�S���5G��K��<{'-(�	�FE4�M{Q桫�ƺ�
O'��4�]:O�����u��O]|�^]�/# >��@��d���;H/N�m.qǧn��	�}�$x0%Sw&�1ߔB� ������-��/n֮ ���P�+tN��6���B�G|�8y���%��Gf�۷�D��!�~�2-V9�U3�ҥ�a�M���[�XA�]j�� ��<�=�������J���4�#,Y^��7^mY��R�a{Փ��\E�(��E۱]�wx�U��e�b�9,=��8�[&��u	�Ѝ�(M����:��J:vR)���Q�<���'#�S���R���o�:���s�.S&���H�%��Qz4`��	XM��x�u�;ƨ�25J^�|�΍��΄�k+p���ê��#��b�.1�[.��J��`�L:���%�9O����
M�$�6�TA4L�|�^-���6����^�vΤ��.�`ֻ��4���~�h�3⯟^���v�kI�_h�f[���s(��R���m�S.ʹw��E&$+�~T��/?C�C�3�fc���	��B����×�sx��jC}��M�&�����ˀ[[~���	�[�U�LSYBv:?��+�*�E㺊Ux0X�cu�x���D�����k�[��l�{���g7mM��4���P��e����O< �8;��hy�M
D[�e���4�)��K��?�x��ZT,\�c?h��'�+k=���j^H�ϸ�X����B�k�}�2���Qz���Xi�/*]�h�r��GA�-��'z�L�\�����Ͱa*c M����;�_ �D�dd$So~ٯ&��
�T�e��6a��s��4S�D��[;(������ƈ��p�{���P�Տ���'��^A�WBa�#[�+�`3���>�A�@�d'!��S�:;=�I�J�C3�u�k>���*���M����_��y���>(&�g��aH�.�@�rk^B)}+�Z��m�z��v�`)�2�J̀ ��I<��ɇ�o	ڷ����X~���!��tt4�2�Q��$?*]�z	�a��ѓ��N��\�JC�T5�W��v֝������ټ���(r�?L�e��(#��i�v�X���J�����BX�<�ۊJ2�O0��#�� �y���@*�R�u�TY��|.$Oy9"�֯*%]Цo��`m�ղ��&��<�@��q�HL�I�[��� [��~S@a��x����5,�e龌���d��-s�zwӕP��'�h憉MO��<�5L	MG{S2��L{�Go3{vܺ#ER�T�Az-E�!�k:�փ,������$��˫m�K���<9�C7:c�6�
0~�ԣ�^?.g��)��O�o!�$�5c��y��LNX� �r� nc4kTLWhp�	�O�$,��7F�<��C�3~��ۈ�$M�\�� .��4(WTe.���?��U�jc@S/<`�(��zڭ[��ş������!jF��7T��*�U���?����?�v����2�:��B���l����Ci�f������s�=����`�8Y_*��v�yg�	m�Qt���yc��1�P8�����`��[�{<z�2@�e6�7�=�\<���B`�G+	)/DKȵl�]q��Ϋ/��Zwu%⪉���XCw�S�M�B��`�^�<��bD�k+=��ub߁�j�R�d~����o"������]oi�Q�P��Y�����{�CZ�p�hC�Md!K��y���U&���m(�h�L�5O��.�a��m���,X�
�V�.a��3\��CR��Jh�Ч2�*'�R]�S��d��tZ�z����I5䏚�v}�$u��u1��L��'BOx$���h�L�
��眖�C@u��i��,f�1L�S�8���5��З�a������w�!`k�l�p�v��
��paU�����C�� �FM�7�"Y�]R���d����$�Ϸ4�(ܸF�Ք|�VX�ٽDN���{4�o;�
,ċ�!�X �q���cBg�Q�,*�$�P�>��H&EA��"d�pQ^s�\�"J}6ƾ#�{����d?h�$`w����yڰU�t���H��ۺF���y	�������G�hG ��u�����2̬�Q��C���>��$Z�C���g}�ptU���5-(U�ϳ%���!� #.��8ߨd>aZr��3�5�-,h��j;r��X`\:�����응�ΕI���������-�#�Vc[	Ѯ��+�p��/Al �`�' C�׻0BB�|HL�D%�+]�ؐ1���Rς�5�	�ݹ��>=�ڟ*�%�%S@�SL�E(��=�r0��R��s���#���H�8 V9\� R�����p�R����_���0������Ҋ|�ϟ�h��zv��>��>��ą�-� 0��.*�k�K�p塪����@�z�e������f����U��]/G%cJ��p���w����,Q�~���T�q����v���(���̄��>8�8�I��|���W�';��k����S�:��\��W���&jK";A/ '��o�U�M^�V¼��C�Z���N�~(7�|P�={�!tmC��'d0������Sdá}�&;4vR2c�=A4tmAm����e�(BL�ܚ�����j}��͗���n]��}�M�ij~��`�j��ke��>&:�_��P� �ݎcY�&!z@� ntF/4��.U[Y�͒g�Zȹ�eZu����[���
������wnbVy�/��AfE�
qZ0V�@�����5�]�ٷ�?�|�v�.�q�K$ y�}�rq����c��qן1��G|�{���Zɋ�奻/�0<��s ��c���KH�C�O�O��`��Q�}�̐t�X���#�&DB_C3$Bk&E�{P�*Nar|�ʢњĹ����PJ}��N��Y����=�6L]�ew����S����R[��#{�$O��$.[�H�3���־'s����Lz�Q��eд����
�50)�h4E��R�54Pr%�����p�y�[����e���C�n�lӡ<�GR%��_Xd!���сW��xfcR�1�L�*_�]L�'�[��å�/����\6��.A��^�.�d1�Wyq��g	���9����1R4[�z�\<�������N�]�T|V
5h�3�eÏm����<^�� ˝D.N��巼$��#�H-�22r\�x#����H�&K~}�YNZT��ƈu�}Q	�gr�D"� �w�cu�>jn���ġ/m�l�s7)-�pZ?�%3�N݆ܚ���.f ��v|h�{�"�#j������Qi��<᮶�0���ا/6���{kA�6ڧ�B��8�|Osg�F�&�S�ն����Ǹk5>�c�k��,^Q���fX=���ƞ�]d�D߆<�[�w��:����]~�P�v:u��\�B��ӆs�%X�Y�2��pfC���َ`r%_���Ǭ8���x �P/~�4Q�+��;�y�y��uT�*p�
/}�l)�x�����}���؀�֟]e��X�3�!uu���v��A"*����?d�*L�ޯ��k��ߥY�K��Μj.���_��T6cp�^��D�E�S�>ߛ5�M&?m����7Ά1ĆU�4�&�m@�g>J0q��R���[[�F���P�x���D����+������B�2~�]F��Ew��hV8D�ha[���\�)����Щ�t8S��D��$�XU\o�/@?q�SLթ�[��:�t �=������3���>0Һ�dr`�D��mUې�p��� �c2~!�s��L^�E;�e�aM�{�{�Q[��5j�wG��Ε������S�R���0sP�@{.��GE�A�J��� Gy$f���i,��j�[�c胓oS�q��[��4�R�Ƿ�1R�<$��`\�����c��\c�Q��0GBH��,轏T������W���<�]�x���㘐H�V��w�K�C=TOfI�6�2 X�3	����\�h܇9�.� �q�;����3�#1q��0�v�,S��܏N˨���SM�H��@�y���N_�]�H"�t�f�Ɲ@	M�2�<`�U$�ȸ�r�1�����ȑ��vqn������l�$⯒�D�%��V�֛��1�\�K�=�� <�@)e�q+i��k7C9>��x������h���3��+�djZAXoӅ@�tU��(�evZ[�w���#4U��� �8/�n�
"��
�ҨKc�/(�'x����P���0�� �X�E]��{Q�B�8�gS�]P�>dX]����zd�sx|��h~)���g�A�N�n�U6���z˽��ޮCT�i|��4������ZiۤW��d����R��r��w����G�O�%����b�J��	����E���Y"�8���e�Ill��z�=�6���@�W��	Թ��Ǯ���V"��o��`�V�R'��L.��,ձ���&�B�0`-Ć5�1OUN����Gۉ�.
���������	TP�r�&�e�%xV\���'"� "��<&�~�k[�猟�.:�E� KɃ1��K�w�d ��7��O
`�������g#���e[+���E�m����Os�>�|�)� Q����m:���?�_#�Q��Fi j#��o�>ڦ�$'���WSwfbJ�m����ufpd��t�|IWn�P�f��������<��U�-��R�~ +��p�S(��>���I�2�7�M4U�TwbŽ:#����@�r��T
���h#�0ϳ�;����l[�U.j���;3��އ7�o�/:�ܹ%|?8��k��^ϰ�U�r�Ч����lVkp7�n'�5it#�j��4&^>D�z�5`)�|� 4t?��(�c��r���4Y�Y�5\���i��8+�4b����o�";�/����ը4�\���+��U�<}5�"y�z|;�"�W����!�K�d�[�<�~�2�֨�N���BN��)�&��P�����ۦN���ߖ� �%|@S�,<��Z_XWG���}ܩ��V� �*�Xj.���g���������h-�K|=�(���4��b=�r	hɍ��~4,��UG���6��[�y��-���b��!���(����\KT;]�.&Q����r�e��� .D�de��!�2Qș����R�2�O��f��?�<9�DmSq7s���'k{��wg'o\��������4������&�wuؚ|G�5�t���p=��E�������͟�ųֽ�K{9.�/�@y!Q58�j�$�}I�F �~)�P��sgLV!$
�e$�])D����m��f�a��N��>��{1����p��)³vc�o����'ם�=�-|�hf�("R�Б��]�N*!~?[�i|0��k��$��b{�������<
��j��b�<�Ϋf��4�c'��o�	�$�:��Ug�mv��K4�b�Px���:��G��M�MH���1ѷ�Le�NX���*�%�""�۽B��Ah�m�ۘ�dq�Ɠ��2[:j,gb)V�ȃbH��6�׼��c��YC��B� y%
��ذ�z`(n���Z�b��e:�PތX�J�ރ�V8�����-�e�>���g�Ԇ7�Pv2��_PC�}�މU�&�6��H��q���[�ʄ���܊�I\�9W�!^t�?qY�1hScvO>dN��D������� �Y��@R���vj��H4�i��Ž��M�MI�%��:n�x�[�K��$Z�g^u��.@�lC��ע!�;��y�$�ͺ�M�Y�T���"�tF��De���GLq��o/nZ@K����A�8<p]��>"����U�*��Y�ߒ)WvQS�*;%��8���p�ޓ�jx���r������T����4��0��$�PωW�^S��v���cd��������80HE���5��&�V.���]胵�˝k�o�w�a�C���7�s�5��{�ן�ѩ�P��Z�#����ƶ������8��u�u������U�
��tFNJe0mn�j��� `�YH"E�J@�f�S�J��e|���rפv^9���s5�[i|,�i�7��|���L�͝;�Zu�[�����1"cD���]�oWQ(�Ƹ���YD1ƹ-\�\�j�E)�i���D��UJ{�9��������4cy������G�V��J�%!�+Ia����&���Y��T�#LM�[����@���H�*�NMk��zb����B��`Y9Y�j��S)��>�َ�pNS�ⲯ�����.�Z�﬘p���\]�Rp���v+ZM��4�RYDP�v��p>@SW�u!E��~t���M痠���H3�g���0]%ڄ8K�N��o|J	f	^[OsZAцS�t��!^?N�_���c��ֺ�G�g)6��$�Z����Eξ��m������o�H�I\�����I�iZJ,\�]��E��Ao=^T���zĩ���+m���t��?;��6h)��~�����v��e��,L� 9��&�W?�+��ߢ::��<�I��ºDPc�t��5��D�8�#`u��2#��T�y�(��>$x��6Qxj{���$N���T����Hd��/����˧L]�#�
�ɌՁ�̾Y44qH���[݄=��+�m��e��_"�ʜː/��"E�1��g��`�-���_���v�� C['+s]��d�xC��Lg7P/��U���C5���Q8�Bu�ص>(��j�tß��G�A׬���M3lgW���.8�1q������h*D�oc� `��sbP1�8n�=�_�1)�������Q�Q_f���F���>�����(�$&��-Il�8��*�m���jUv�-��<��튝:v�	�򌷖��\�!$F����$~��\9	;�1
J����^��o�<eaԅG�aFQ0��6\=��?���#�����O�VW:��� ��f�'�ߎ
��|I�CN���U��O&���7%a��T��fؘ�2.�͢ G��5���e��7�~��I�{��;�\�N��v+0�Lh)�u�Gwɱ�ia�k����E��}}�8-��m+�@�{�+��&��������]�������Ҍ[5_�WK`4��) 9\0Zx�b�n(�b����8��&����9%���"�~$�K�����K��,p͊�"ܨ��|Q=�=6Å�l��$��;���F��Cȼ�V�Q�w��{D��1�n=EvNgU1%�^ ���,��YH�[���f
mR�y�0��Ż�I�X�J� >�6��X�U~�:Oq�ʩ�
~��*W�1*C��t�g�t�
��2��R�0ʁ�F�裲Bs�	�t�X8�,ԃ���kG�WǞ)�Q���7���By�{��(/�r�8���G�s��:	o�H��͝�ܘ4Jʾ�1���"�.!�U��.r�}o�gU_O�B���I�s�GB��.t�f��t�E�ݠZB�-���縂���߿v�C�K������z����y���D ���d��&?�Αu�����_rc�$H����ͯ5i�����݄C[V�/9q]Iɺ:�U�QJ�R��7*��=�BQ_�e'Q�ۑ���� �%���u:"·�n�K�Ey�{}m�+�kXAq��ɭ-8A�(�#g�S�#�ߗ
�<�f^@;T�r��Ƶ(��eی��VS�ԊgA�zM��-�B��hj��;DTnn%��fdL4/����q����iqo3�tuTB����o���>z�'q�����SH�6�_x�xPR"�M�|�A�&k���N�%B!R����i>>T+7�֟��lދv�Q��_�G�q���D�S%bU��	u*��aϖ�����z����V^ ���Ć��C$I�G�Vp�wy��!�j|}v���W�Zxߗ˜�ٴ�\k�i }q�|�7I ��7#Y�V��\s<��Ow���6�V�j�)�Řdx�|�y���?��+�Um/�ȯ�æ}��ܓ��^>^�XR����O��Ogq���"�B�M�q��FrJ `mc����|�����r�H�ے�W 6�|2zS�*aY]�̞�ANi؝��	�a���s�8n���-ǒ�*Q��A����t�?Gcpa�R
KN�X���?:.��}�fQJ/�
�{
�y�����w��j�3ǎ��qs�=����`��1��&�au��%��8�IK�����f�7�$�W\?�	�����ף�d):q�\�6d�rj��'��R$Y=Y>GR��0���!S���G�.1�B��(�(dЎ�����AX����Rp렓�}BG�D6�j3d�:ch�{��t�Ve�������$d�׳M@�k�����D!�*[G��� ]=z��f�3��<>��2el��[��ی�� �~�B�7�.���[���N��9l�����m�F��4�5%�z�P��u�G � ���LI�*�+�QB���T�����}����7cɔ�y���`/�7� ����8��N�lld�(����|���g��"�����q�zK�s,/�����/�&�Q2�@�T#��q���?�c9��.`Y��w�ɍ�/k��0�,�l�ϽK����K��0P��bAj5�:�r}�}���*�qcN�S�� �����5e����S���3��5�[a�k����V��s�.����z�щ]gg��L=w��V�.�X��.>�K�aK�J���`ǥ��0��e�h�w�)1�	���o�j��n��h3U�x�N��B�O��C�D.��� ��+zۢ_�H9L���j�qj����E&����ʝyv�;!9��	|w[;ī��
�G��q��f\�k��Q�XBf�~:m�\�/�^C{�~�L�d�6}TW%���I�U5�`
��6u��'6�u����0�e�n���}���AJGU�W���wm%A�%E
 �h-߳I���F;|��䔆��C&b��s>s�潣����ޏ���È^��Eˡq�H�ؗ=�UӲ!n����@�J=@�~�7a�J����pɯ)��߆Ҧ���Pso3f��H�<�+ɚ�J�ﰳ<,�0v�_��c��2��ό�7h��j��k��F�WS���W�;u�O�Ц*��G�������>���Ｑq\�B���j�ax�&G���~*�Ut�[N��.�yR�¦S�����4�U�nq����}�W=X��n0��Үf���X���y���>���|�ߒ4F��De�d��i�}|�#!�M;ȍ:r�||��╔�Ry6�TP�{�u�1����wH,�F/s�|�|W�l�����*x����9D��g�7sG�j�mu}��r�ʣqGA�C������LI��p5�<�{��῝��S���i��\�s�8M�6M��[���2�Y���!�����db�M=?E8}�6�,�A�G�mErz�3�K}�Te��}��P"3/L� �T0{�~�D���!	>��a��3�b�"ο%�Zɘ@pV�u����lb{};#����g��`)���}��T�|(1�1!��D	�(��Ά2���#]��7��u�gjS\�i_������sߵ��tĩ"�y���'O>S<�ۢ�U�=�Ω���j�䬣�����*OI�{ڀӽ{�~%!�W+!��)��l���Ǐe�qP~����QC��K��(eM���9��	�͢��H����GY!{�r�pma�5�(I~�撏�;��fgp,�Yx�%k�nf�3����j����[v:n��O0
r0)���Iʀ)�a/T��-G�fΜ�֐���Ծ��[�����ف�",�/s5�5�8�Hcނ@:�$��Ѕ{�lM>�x9�������;��7��C!�x�DY�c�����Xg�������~r5|'F9����Ԃ5;m=k~�8{D�	� Z����Um��U#���O@�˫t��E���윻iP�˼���W�s���8��/�a;7�
M�x��I�ܥ�� b�wp9�G/8��˼�{wy���U=��|wa�mq��|��q�J:_hE��|���B12���ܶߜ���Ϳ���iW� ��6��i���}�F��G�g��o���{i�n�5�T��}��\�[�z{]�1|p�鵎P9ʰw��TT:g��RQ����0xZ�+�Qp�Y���,�2:��ɱ_��~,Mfjg�B�ELl62a&6��$��
���9��+`�)�է��-t��ơ��Ҏv��2w��z�x�
���*�(��L>�!����׵��?���մ�6�'��{���������l��n�C�V�z�#���C���}��<�m�\`�B�N����=�L�e� �c��7+�r �k��ʺK'����a&41v�����n�|��[�R�"��T��XJ��0����c��:�v-�����j���6��!����	 ��%ٔ���om	d�-�㆐;��T�����(� J� ��x�JɮUh�$Sv�i��U-���)�e�81���*�^��jt��1����G�r�f6�0%#N�%H��f���ą˶������N��	'gBQ�z��� 1��ռ�鮀�:f3 �N�����I ��hZ9ٔ��d�G�V�,��¿�XG�@�ܮY�b!��1ӃsJQ^я�2�{��ols����G��e�����ģ�}%��o�����z��E��͇�ğP�{�	�>H'�1|u[cBEw���Ү��5�K �Y��.���7`�:��Z��d�ueY"������-�������4X�u%����m�g~�
)��z`cr܃K��9�c���J�k��P@���x	�ۍ�A��k��Rd�ֱo��tS��64�z��b����x�W{]3��h�u���.����k_����t�����nZ�' ��pB�*�%Q���K��dS�EW��(-F���%�v�U��h�K���q�c��7T�)�g���yNf�l�ܾe��4�/�퐀����{���#yud�}w�J~����w�^�;��ý��i`�\�!��2����H��gLHv�������d�k�b7�+k����2���QM� ����;u���d�ۭɎ�\:m�ܗe=�^�k���� !�1^T��t,�S�|�C_[��R��
GY��!wχCۨ�j���w�4E��d��x�a�0���)#�u�(VF�hE�!-	����U�A��s�#�
��f I��^��^��M�3�dn<	2�k4���"t	?9�
��rUS���8Qm(`Y�����m��GK|��\��V$dfo��"bT{��J��$=���Ȩ5�l����d�⢘��qI�:���.�0��܃ٳ������}5ѣ�bm��Ao��i�®5�A�cpL���-as�1�)t�g>�/ݹIUVueY��T�ꐳ�/��*by���r�MO$���}��П���Wrȧ���uYxl�N]��FʑF¶h8��vU��)K�K�=y��"�Z��O�2T@e��<�@�����Fbo3�U���6��u{�/&��e�p���g��>v��6:I��@�B��C0����T44�x�̖uS*�2�.��� (ӑ�3�踌�zR�v�FL�,D��K�}J�l0o<)p�VԢQ#�sϕh�HE�~����ʺqx4���Tk)���::�2���҅x�rd����>,����_к�.�{�ۢN��A�_���烤���4�Di�^��C� ��렟	1B7<���2�s����2�cՋf釄�=�?���,�o���.��uS�=����y�~�D'b�<�	S��RGG�^��U\vi��8��r���P�k@l���!�Yw�~lǱU6"����� X~�unn� �%�2�8�R�DTz��w�d R�G�<x<xI�U��9�n�Lڼ��8?�!�C�O�6�b�gF�?���^��@@l��v�)�}^�ro� ��}�0G�OF�~�{����_�,:;�j�
d��A����<9��rG^R~"�2>X�c���F�Pl���a[�C�ű>�S��b����(��*H�X�-�,�ד��]d�mw+�6��.��f�5�x3�^�Z�zn����wȹlnr.�S3o�T$d9(QAɫGO�<�.���x�o[?(��`�0��VRO`�ʯ+O���~a*)%X��20�&�vc�~EJi,)��F��&���N�	�w�x6f1#D�X��D��|��r�1whʰ�t��(@h�1�U-uA������Os3�����xGC+��~��Aͥp��[�}��}� ��5��յ�SO��+�+:��u����;Nd�sw1%�6tA>��ۛlɇu��J�����!�V�çǚx4�͏�,�MRL���|����������ꘗp���b�4�>V�9a��\�m�v��8v[�c��w�2�����}�Jb��7��ʤu�������6��A�/��%��͞�?.M�S�^}���9��m�YФ3�ӯ�?D���/o[$٢3�ג��j��ji{3m�d,KvJ׫��o}��l�\E�?_�����0���6=ir�}�B<����*gro�\ŋN�1�`��S1;tn�Gje��f�B�s�d��ls-k��D-P4
��d�^adR>Iw�-�?	��;��M�h�θ��E���y|�SB��E�j�d�U5@+e�<�V�y}Ăj�a�^]�s�Q%�WEa��r�4NV?H�V�Ec9�7��u�s�-Hu��`�M��pFLE�䎷��P+.d"�Ϲ�\��7����BY��.����M�z�r"<A��K�}[>n��3q�DEI_W�
�T44��ug�����Dz�?5ʪďA,��B)��H��Bؔ�xL|Z��<4Jh��NH3�WIu�+G�F�G4�؝�5��{���wA�v�0��e��A%�k�~���/>�[�.�L���IC�15�$�=czI9�𷙞��|if���?��,T8��7Z�:̭:���:"�z0P��;�S��F��pF�[��~G&�VD�e���a���/���{�ͭ#Q��y0k�	�ǣ-��Y)� ~����0B�-G,lQ�҅K����c�>��|��9��,R��ť�?@�S{��?����m�Lf��FC�?a*�1a�XC/޻��" I�!4(��1��i!a�$J��i �}��>��}��4[��V�`��Ud8E[�ym��X�&�s��@Y0�*ބ����x����(��?���k�w	h^ϡ��!�`8i����g�@���7A�+�!�Jn;�M��$�٠}���s����f
1:�2�Τg�*���R��Cd��K�SW/	Zm�
��7P��f�%�9Pt��v<<�c"�1�d~0m:[R�A>;��x��fꟛsұ&�=|����+�6+��G�i�m[#Y��f=�[֊}�-K��������>U��jhIH�+���-�e!]>&*ʷ( C�t�+�h
��q�@�~��� ��(���z�ef�߄��qO�?�;meܛ��M��'�/��)�H�Gf7C&��D��1#"�X�h�f��1z��ΒjǞ��Y)�8t�ω�#_��춚����tS�?�B��YB-�>:�qr;4&�G�����BW�����p���Y@@MNәM2Q��O(�9�ć�C�\��oXI�C���9�`hM�l ��U�^<�t�wߍW�̰2+�b��sc��p?�Bo*����Z�fA��{<d�=��&'�v��I0�QѾء6����ޜ�����e�\��9�@���َ����$��Y��P��/�"�y�H�ځ��K���p��@:BW���� ����-A`�8���B�@Y�pr��,GE�;�I�韁;!��{{�@�� ��N��'� ��*Ҵj{Ž��`�������՟*�'�ю>0B'P�z��E�����<0ݡ���e����˷dz�"�a�;���jD�L��=GM�.��¾�����1�pЗ�km"� ��׹of��T���W*4w�!G��)ж��)Ϋ�Ð$�S�hZ�Ԅ�!`Y��S϶�@����5e�p�!��)��p��"!a'fBo��URN�k?ƧdZ�Vy˿5}^�M����.<y��J��$���&l2������$_D�;�Z ��5����ϣ�����
/h{��~��G�?�F'�7��y�N���i�7����ᣣfOG��N������.���f�p�5���c��Ex� ��&��V^����@����U�Rnƫ�cb��*�A���+���;:SC;������~�h39��$o�I�F�	l��T�4�Po�U���K��=��\y�M��{����x8	�*藆�y��wǄ A�"�^�}7�^�c$��;�.g&�'��l��
Q�yG[WrUU�L6D�H���&;t���cF:DL��)a�e��U}���N���8�wN1�]dR���2)��ds׺�z0���7���J�+h��~͛y��"�B[����RQ��f���IU"��1�۟�'b�ڠ�*7��oϽPP���l�uE�I�U�\�0�����=P���uֆ�C�c���`�|��[��-d)i:mJ8�]�O.J��tE�"��і��M�&���I�,kAId	

��Lb��0{��z��8��d�,��� �����qU�Ř%�z+��q�-�4^��ˈ�Bh�Į�a1q*�����W��!�w�|����_��7M�tO~v�	"b?o|	�\��Ľ!�d��x@e^�N�4������?F;_�yk���%�CLk�6���h�l���]�O�+貁���Lв��P��`(��/������~�����Co�ϲ�pA)p�>ؗ_ޣt)=	5⃋߆�rNU�s"{X�G�˲+5����Ʉ8���m��)�O�������U�S���?�g?u��eJ@*�?�!�6�P�ȓ�u;���A�O��<�!�l�9���69�v��N�E�����]�W����gs3[F�o��:<�
�]���V�����2��xJ� #\��qm��pD,U�3Y���j��~IZ�M�Zl�����bN
qw:P9��k�'�GJpQ�[�e���^���� ?��)��C�.6#��U��ǌY�.�C��N��E*$ü�% ���$�rG��fu@��|i3�G!�(�$�2�tF�U�@��p\�Vy�����n�-��z��DN�@p�̑��ͦ"Б�G��w���3�ݾ�bֻeHz��o[@>a���S���P���D!x�φ�* p�Z4�%���w��&��G���	q�6$�tw,^#���_��	�����]'}�������E/?d�t^��\���U,fQ�غLZG��;i�Xedn���8J5���@T5���!�J��RSo�D�+Yy��B��_I�K�t8P�O����)9��NR1ʵ�[FUt�;�~WCI,����@Jy(�#�,ыh��;��R.Nъ*��	Xt �\X��
�� � :e�aq+���AsӳB}��A(I�L{��<���*J�E�SJE�2w*6>�yC�܅b���ݑ��=�,7c�]A_��`�<�doF����Vl܊�ʪw�@��T,�H3�m�0���gt���Ys���̖�}�T뉨A�.EN�S�g��b4�@��~L�]���?;�6���N�*���\@r\��H��ȫk�ߢ�p���h�7$�"kg(%��ndh��_{9"��g���$�~�^���-���!֖i��b��y�{��n*(t��6��+Vw�(��R~�_�Ƣ̜��^g9�M�4x����4�)/#g��\��}�%�Q���(�������ܰ��߁,y�v�L�� .1~m�d��L����tB��ϩ�3�D�fH��,�]�8��.ŏ�X�'�圗�g�H����������b}~�R�ON��X}m�u8���Dn�Q�y������ 蟌�kni
5��Į�h[DĆ�0�M,A�l.���fjAP9�ꚵ�~�|d�^���v@&�t"�w��� &���Y���Ќ�~��u����n�x�A����e�Y�ʸjlF�ly2f��<�yo;?��p̾r{��p꒼ҐF3H��GP�m~t�u�*#Q`)�?����!�K���)���b[�.%��H�9���y6ywO��tǠ]��U�_��w�ί3�x
}�a�̊-�t�� u��u?��Iyf�����q��=�i�~sۍ�����%n� n=�+<��>��-��<7�st���c����@WZ�`L��;Q�G$|Z	���@:���������.���C>��yʙ���!s�NNi5���*Y���k���Ǉ�@>��E�wu$��i�M�fP���2�r�NޠV�z�)?ӟ\�b��L,]�n��Z׃�Th�\��QBnK��Lؚ��<�ת��U@~)�&�`]8�?�������u���;�l�u
�J�≮9sV0��5�Ll�Z^m�F��)pw��*&Lā��גҿ��_/��c����:�;Fs���飩��l�ܢR2���b���o�%��fٜ��0uA��8��-��B�=#ϙ�̪��1��\C�l���x��h(Kւޕ�o�'_�ĖyU�VE��l��Ύ����>�}�J�o	V`��a�k��ɧ�d4e4Y�LӁ"���G��ѻ0��wgycK6:�����7� ������u��}&	+c=���m(0*�Ow�@�*�5�i������.Z'Y�|SB7,���;�D8|`�	�W����m� ���e�ݰ5�� =&��"u2t�RF�5q��C��﹜��a�[�+˫�L�X2SkVk��Sc�����`$��#�< �$aᱜ$�]E���%��?�s�7��������� .�ؑV0K�=7�2N(����W�')���R.Q�f����=1ܩ<B;@�L����LF�/�W��]���˻�y��ݥ�t��<*���헩�aN� 2��4���HAeȪ� �d8�Y�"G_�`��:����������@��
��/6�:ktL��]�Aou�������O=��X_��F��:�?������AL�a�ٹMq�� /�O'�|����e=9�P�j-���e��T#��p�m�L[��ql��|��b��+�졉�l}�k$� `d��ݝ�w����p��a��L4@��o��?��:�#�3�)���Pyo��o��UC9�e�`Y��1���Ͳ�)vL���!��C�y\��!���@�]��H^~0�5��yw�=��1�O[��{�p�^
A���Y�w�?�ʁq�}����h�mt���]�h).h�<�6��s�D��� ��}�]iܾ�YA�V��}���q_��\'�wv��` s�@���%�kca܇�kFB%Swb_>�`�n�f٠��$[
����oj��av"�`���F@����� ��d����	�������O� w�ߥ��*�$��Si�
{O�y�%&���Mv�T%��{�����fw����g��P>qj��V��d��h�f�;O+�6��j�F�pNP�t2
i}d^D�(_%���ۨ�j�t�B��� .'|I	�rCM��Jo�V��5'ꠈ�����>�n$v�*�xI�?*����:\�
�5 a�C_�&��q����d�`�׍�7��E��Pvj����q���ܰ���[�]J@�:$|^tGO&�hJ_��V��SG�r�{d
6̨"�K\������(��=�ԓ�f	k�������d~<⠮M-���	�5�8�\Vͽp�U�ڤ?�����P0��|kz����sb��x���ltz��j� ��R�թ�N,�}��]�s��S9k%R\}��ņ[K�ٚ�T�bB|T���l���/S����8-��	�^��	�������[�Z`P��pҒ����v��S&�A��A�vd�؅��3�����um���9B��>����
��jʊӲ�m]F���<0�����u4�X�@��dc�pgf�M{���I��c��:��k�������ΓW�#��#��(��߰��g�v7v����.����u�U��wꝻ�WN�3t"b����LYW_ L�oi����K0�����dFtS:+Aܻ2'v�_��Qe䢬���F�y�zhC������P|?VT�)lp^���2]�0*����=�˄�BF�߰��D�Y����Pn�^tPk�&y.�ƃ[@��*��hݤ �
�Y9Jz�5���67Z�5�F�\��ZZWSH�F�|-.*&��h{��B8ykόQk����Ÿ�1�٤�r�;o���L��z�5`�t\��?���)Mo
��1�A��&�f	�P��sx�7d��q�0��&^�,�Mg��p������~��:C�l�he}�(�g ÌMѓ�S�-�e�>W;�Jܰ���8��Dv�:G��O�!��=�?s�-���*�kG��I��-�`�Q$�Y峳.-*߭Z�,��sA�Vޢ��G�B��5��̑з��#��ņ��ф���)K�� �!��̖��(�}�YJ^Ut�'��mQ�G��I�5s�`��~��O?�}2_d�>]������`�ɵt˭�9��}j���}]���6w s$S/Vd��u�0I����ae���c��Zy����oW��@Z��pÞV�Fr��ʬL/>s�-KG2ߎ���9R� ��a�׎�uժ�W���z�r���3&�fdl��"�l���[�S�q��Ë����ioL�k<�!����p?�hR��A}kF>XB��5-������'ر5��״�16C9?����*���:��L��͚y�s���:�2��yl����n1n(��ՠϕ'�fu�#�tiF���\�3c<kO�� &#!:�$�J���}�D(nf�~��-��GDfP��K�I�nv��zy���)�}��Hv�4W]P�z<������Wγ�bHr��-+��V��~�ӄ	>=�j��#�-��ˏ߆<ɛ!v��w����yHm�acb�t�U�=�"�g8" ��و����r�n��g3t;JBMf��L���Ъ��N���^�ի����_���qޓ���e����ե~�c�3.�d'�-^�ų��cboT�M}�1
���8ƃL��0|�tT�����l�e~�_�}�p�J>S��V�E\J�/T,�{y��~���@S��f`'�=��0��ix}��&6QT�z�X�JVc����dۈ��ق>���އt�B͉�m��7�R��U1y�@x{���!Y��7Y�l$jUa�(F�*-o�����;����u��D��]rVОNu�Bp�:���T'R$/B��W<u?w0 ���YU1,���w+�����\z��˨T2��5��yKq솚����Mi�"6v��\�SQgES�/T+��������{OeD\��m-ɮUM @#tCv�58]B u���Qr3�b�\�b7x�b&��N�_���#.�.�5��p��m��f�L�҈P�R��^�c����@��ܩ�$�d$b�m��v��`y�o�����/���D�6h���jg���Yg�Ս>K���[n��~p`���B,O� q�c�@�j��[��è) ���9�ϔ�Y���)f�ܹ�������b�κO�@t����k
��1��1�&�f���&��̛�S��yn��� ��.�����P��_���;����ܭ��y��B������D�Z�L;T�c�ޖ-�% ^2�g�9�����)���L�磂'��,1R��s8B�u��3��=��˻ ϫ�ӤɒÊ)�2͝Z_28��&1Ί\	}��1�G��s5��Z�.�g����.���������f�&hR,ja��"��4�#ɽ���;��9�@�,	�ç�J3���?(�LB+Rܡ)��X�s��oY�O���B��mv��3�����Wyc$d�N�+9�{��v�/�X,�m(�D��xC�t�fx�Q9PM�^���n�Y4!;��ԍj3�r����%�S��
��Z�^�4j���afSAa�hy��Aߝ��{F��1��^�sv��4ؼ�N�����}s�6uS��\'�Hr�D��&��m�6T�6C�(
�
�+�7g�N fU�=?<�y�>�\$�ȅ?�0y�n��#�	k�Py�+ɵ�x�9��#t�1@�;E��<�ڑ��蝢�^��	�,�^g�g�R��w;���=�u��)0�����`��ޜ�Y닧�&y�x N!�j��v�S=~��׀�0J�����8.�S#���gљf�?N��KU��p~)�u�vL�����{�Z\ѻw�V����pó��>�b�����S���)vz�4�q�i76�ʾ[Kȉ��:���,&���'�@%`䙨��]�v�j�ᗭqф�k}�Η�P�-�b�m�;�G=/#�C���2�*����'?��R'%���Jm�n��/{��P���Ȿ2��\^+�Q������[9��"1�ћFΞ�vl���F��2�VJ *�!K��3�Z��;����~�۳���9�$r���T���A�'8��k=O�Y.4r��4�>hKg�\�H���L�p�~<�p�L���Do�[�B5I|"PH\%�W�-�'�*Jn��=�1d�e��эw�rm��	���.9}l �����N��|jU�aQ���it�
�������*��r��٠��̛t��U�o�kӔ*���6� �J�s���bGp:.�xgD�G�|�$�	bT;qf &W|�b4��^ŀ!j!�i�e�i�?W*��� ���'�].
��REƊ�=e[# ��Xs|͚8T��{�����ϹW���MӼ��Ԯ�e�#�(�j#x��f����E�Q�-�EU����g-G=�U�O�D$κ=2�C�!�[V��/*�](fF�l%	�W_h� �BKw��vB��fR{~��O�\(�I�ޢ�=Pn�-�T���ˡ'����1����l�<)_c�`Ρ�<�R2�����R����ݼ��Kk��Սi4b�!���]��飥��8F��Y[70%2��9�X��~MV�?)��>(�:m*A�Eu�H$Ǣ�U�����܃Y�F덈!����*�i[�ݦ��[t�>C��9�Q�ŇFއ瞿����Ը�
�t�'�ۣ��p�d��\멢ɟ����Ơ�� ��1]h�S��:	�R�Y�� �ϲ' L��r#o���8�7�t���c[fx �~u��ӅC5k\��xj��g�SE^hߖ� �����������0�#�Qr�u�Ð9,Ҟ���5���g)�څ�x��8�VK1�X�h:"���6O�d�'�T#h�9d����|~72E!�FPտآ���3&@��6�Ū����z�E]^�~*����KɃm^{-��e�R�7I�� I�w2�2���3���E�*4be<Jd#��$��O.ʳ��h� �d�zi�#���VG�@1�	��(	�I�ڠ�6E5���n�l��g6���4�F����A��%��dN\i�㨮�Bq���h#@K
 >(�4��t5 ��}Q��|ި�uD��m�-E�cX���1��YuS"s� ��[^����G�/�!
�U�+� c%e=,�ޅtjQ�Y9�������c�>�}sR_���m�2��f �� ˝���7��r�X�?|Әɧ��F�.��kx 'Z-Q7�,��6ae��'�����bZQ+���Eb����Y���F�T|>�m��Ԍ��&gS�uF�{u
6A��=м���p�f�0jy���sߘ��d��@2�z#x���N�#,���0 ��W v�����RA/�@����B�j
t��*S�@M����W�) �D�3����T�>���<S�;�G¹��'<�=��h9H�3W � �a/ׇ�-�iLQ#���լ�} ���Q�{ס� !��ݮK�[S:���)WI��!��� � 3i�h �֓D(�k�vAj�-�K�X;����긪�tvǒ����+jҩ�X���~�a�o�$�kϋ�H]�?���KP�/��Q#-�^g%�3G3��r�	�5�W��}�d+���G��X���]J4V�� �����X���t��l_Xa3H�X�½���h����C3����p��9ڳ���P'xI=�q���˧! �!,oRs�c]�+GɌ-��
5�!sW��� B39O�_����M}�of��Fx/	�W�U�汵g�!'�,"�|a�Q1�	
��r�s?y��<����?y��y�����c��J��.�u�}$>����1����Gc�)AL4�Rȣe�H���wr��-��n�*%\6N���l�y��S=Y���"��+,�\ 1���|PP��䌞�|M��������ENL�[�d��2n����]QO�|f~gu�W�f��Q���e��F�ρ�B�WV=F N��*��ܱ�trY�V���x-�!������XZV9E	� m]�j������٢n����0�PD��I�Sy��>c����*���A������roh+`q��-�Y�r�!�EGt�|h���!knњ礨�±����'Ng4I�g'X�UO�<�V�- ���}��I_Y������������f������
��Z �n|��U��F���,6K�H��+��2�I@�.$$ı�խ��(�b�����~Ol5�j)T�u�3J1�Y��=m�[I-�d�c!L�y:@�M-�-���`dk��aj]!O��\A�����7��b�b��,"�5}�A=s����Nj\�3���嶪9L��w���}d#����T�ʳ�Hz��$h�Z�Y�ͣM��KX}��$������z7yQp��<��I�O���.x2�5e�+ȕ1W&8oD_���Xy���NЦ�	�%t�̹�s#�F�4��	5I���&�zn�y�!�l2��_vR���������%�9�ݚ�J�i�d0W�J:��n��Ȟ�l�M$�@�3'��1Hd�i���Iir�)�6(�h��W׆hs�ܿ��)�JF�g<��<��~g�qe\�"��;�\S��j_@ʁ�9�K�;$a`q��G� �>g#�k~����v�Ϟ�x�r	 ��r+�$�n��hg�-�?��1~7�_���h���v�9���lv��)y:��n����Sg�bk�Tt��"���9��4�X�j����V�)�
�iU�;���_�e޽���	��iNUxG����Y�~����=���[�$�z<e������@���X��@�t��!�v&�aI`��cL>�"�[dG1K�:�;���ðr�	��UCHR�����Kq�7���Hd���0n4�{԰���� ���F#bg�-�����-�̂!x��S��r,�i�Bu��R�	S�S����( #?OZ٤�V6�+�P��L
"K-�R�\ǝx^w� ��ΓDb���I-�k��#��W��aT�I�Ed&%Gb�c\Z�@t/Ϙ�^�����y�O������V����&K�r��b�VDdbj5V�X���l��y	���=��3����c�oP�����U�j�z��v[c]�_��ܑwy�)V;]���j	)SU���+b|�12j����!���k��$�Kz=�.����١��� �(��ڔYh�cѭB�X�ܪ�}��!/&����E�n���q�!}��p��O��\�'�4���"L^�_����I�,W�Қ*ޘ�'"�/��Fh���ǎx�r���݅�y}4�+���e	>U-�?����*�'���4�'�eHH���k63�IC-m5T�
y�!2%�A�8ȩ�l�J�\}�	����l*�Q�R��"䄀��uنM��hl�M�dF�#;��߀l�j��B��k�KC���)Ą��>Mw}��ݓ�,�W)�O�����*�d˃�>o�g6+(�YYS���=mի��A��$��-�qz�����+shBۆ����#�����o�� X�R����XH��j���V��<Q�� 3�*&q`P���?W�M�z�,HN C�%� �ח�G'É^Q��S��6�ŋVc:ϔ�P��)�ƈ�2;�y��UĴ��'��f���dk8l�i�!�&��{����Xi<`F0�P�b�٬��n!�*�yc(6m���V$���`���Vp}�����cS螁e�ѣU]\���)�O8�آ@�I�ۥ��-g��s�2��
X�ѤIO�K�K�F�6�q6�e����7�5�b�=2��;:uW�"��mh8#�'�n�\"i7i�È�����'��@MOᅳ�³.�p7�{��u�-��8Y'����Gq�+B�p:0��)�
��B�J�X�փ�<�mG���B�V�q~�ؔ�ز��*��g+OS�|
e��w�s���>���EfS�T��/�����oj�_�_�����x�)&OFF��Sfw�q���*� ���z�D����ʭץ�L��S�5{���S��S��z{���I��H�j��sRJ� �I5`��ڑ�;��P��A�;#��=�	o����Y&��8��b���xF����$f
=��Vj��g)]�?���f[v�8�5��t�KI��2AE3���͇�o���A^[_�IL��e�Gd��@��n����ÛM��Ų���ʃ"�U(��7"���0��*�J}�Z���J)�J�ַ��L�Hb1���vw��I5�M��q?J���:w����^�����M���vH�d��<��aS@-xK�o�s�/|���wWϷ,I��I�����-�ĈAW�\��`S'���(F��Ѵ�ºAD��V>�P��椷��l�c�to]�����+�����wp�����>�FW�� i\)��YC@�p4ܚ��]�,R/��Zii��R�	����[�d��P�S�1�b�(�k�BĨ{'�ej��ż�=��ic���b㜪o�a���pU��"\73����/�K�H`�Xb�˪�.�2)j;�ckES��-5]K?�4��}&{C�}z�g�?@O�%��`̤uuOX��V2���g�9
��73�E�s�*��θ[���kBC��ntoV����H'����PJA�UP䔨��5�,X�7iۆ:�L]ft1�ILE>���F$�$I����������z���=���A�;oܔ����#�!C�l�')~�d2��$�.�M$�z2ݪ��l(�ޙ�^��/J�|�1(���ϼ��a2R�H? wb`�#l/~��+�.� M0=w��M�۶�cpcD:޾{�;��X��4���-�t6n�un��ǧ�,*z4��g�j=!�M�:�U����WS7@��5��Zu�C��$D[$���bD�>��th)Q-'��5��2�(�K�a�_y�����޷;f �TD�bB��/�1��5��	����Y*�;ń��˜�F��jU۠~%os�j��n�e8���x�H1�
�f�br&�_�z�c�
�Q9�(g����>R�.�` �X�^sCû���]&�00K�,t9�׫��kyv���SU I��4{*AB5Y �u��FSZ��-�fm�g�/�5n��B�?��25�)TQJ����qPn���!�rgjLy�2#M�oRg��H���pi +`����QJ��u�����8����m�ϸ�I�L�_
9�4GO���׮=I�D���bz+Pa�)���J ��Vq����jx#�I�؆ �F��7�h�W�e�FO�VF�J���L�^� �u��e��(��jHo<�@��?�����|MG�΋B�Wh5��buB(/�@���56�_>�[x����k�-���^u�Ю��}�p�j6�;�a	�t?�ދ ��7����'��t�19��@%��,�����4�ј&OӀ�f��"N�3qH�ΐ|��#a��	��#�������=���a����A�F�f��[��X.�>�
���]»�)0%��i����Q�i��H[ P ˺�TZ�y$��Y���Zp��N�sA�US��K�ψ`D�+}��kT@|J���]���T$��Ѥ{����j�X��kB
*A�5�h�El��b��Kn����O��`g��Zk�O���� d��j9��W�EK� ԧɅ��v67c�����(�dq��.y�JKjs��U�R�:o7h�KS.��wB{o��Lt	�Z��<�`�G]��z�&w��^��wh�������-�d�,lɲ��Mu�Bva�(�O�>K�Z��B��JO`:�(�Y]�b"8N�����BlK��4�B�h��+�k��7˻UR�KB\�֚�o�eu���Uo��z����ġ	�Wd3����S�|rXnd4I^N�H��������mx93J�d�f�b�́�jڂ�ji4|����,Ʉ���sw�hz��e( �w��ˁ>����� �0�ԡ�}c�sذ���,=�k��ij�)��x�s���u� b�d�	1�̂�t|@�
Y�o��gC�|�ǘ����4|�D#E�������� 8 nL7����g�v��0.�����L�xY��J�$� U�B��o*a�>l�^��63���M��߿����q�N��Ę3F-t�^/t���r�r�K��f5u>��J��3�] �06��-7�h�^#uc�:;81	���#ŗL�=¬~��M��j��+錂0�U�	/J#�C`.����F��#�<Qw)[�|@��g_7�+ձ�GJ?��qK�ȥT/�pƬ*G�@���5 %wA����"��N��}� �]9���@`�t�\oRxb�o��v�4Nnk*�,~�&Y�(f �j] ��O��_��}��.ڣr6N��dA�{�+}��]��8k����o}��ZF�u�Yf�� ��2��.�W��н/
�����غc�c���p۔�r�?0Ji����W#'�Z1pGsky��l��*��W�t��Z4l��W:W^9��L���.���G��fXk�c�\�B9�R;��Ěc5@�bs�tj!x�N�����FS��m1\�ȇd�'��e9�Gbj!�-h��?:Λ9���X�Jˡ��n�Y+㪉Y���U4xa��"��nώE�sU�#ڱ>.���s�<�r%���h��
�a�W�/n	T! �փ�:���"���7@C�����W�"���}����P,�r&x�o� �*3��C�e���ىu��B�u>oē,l={�
v���Q	!1!�7FԚ��>բ�D�n�|hkz�a�n<�kb
�����&�yh����
���
]���G�����2�:���#H�t`sтb��i���kovJ��6N�B��^&�X�q�X�+\xᠠs�3^N%ӆp
��{@��tr%e,�P#�Q9k���y�"Tc���H(m��	K(���_�@Hfw�@	)v~[q��x�i1� GI"D����͵���� t�vʙ�B�U1o����^g(_�8��	�*��2�QM�T)�D�qC�������9��v2�XD����X�w���1�Q�#}�Հݫ^1�.���(�6-�B:?�Aa��V�F�qwt56��G-#�C�ˤE_u�eպY���Iu��A�5<�F[p����N�J�"]�t�V:9��$�!c>�bg`��}ʍB�ג��:oe������׺Z=�	"��	�Ӝ�&i���':�j���HT뺹�[O���^P�Jf]��];ֻI��p?>�`��}3���C�L^�w�,���M.v#,���b��gO��oB���Y�W�KY�>��U+����l�ăG�F���kh/�8� 8����vgr�fJ�'�B����h���h�H	%#���f�����@R#P>P���U����=-2�����Ѐ�L[�Ի3魑P �����a��b"&��SV����c3�����X9�R�-��z��<*c��]M����:�v��$�>�>�6����B�'�Z�a��R���^��y���^{g~�u4��5c>�2F~�w����e%�'����r ��V Ԏ�}g��]�I���8'�:��r��K�u���*�ԓ�q�ԯ8\��	�IV�����]��|��=��01�(�]��;�L�h�1����8���I|��`��[
�N����$����υ!�y0���r�:ߖ�c3��k|��x��k�\�E""S����cI�IT�m��c����k� �d6�!(����Яv��:ܤ-���;5yQU�$�t��dn�|}��4J2]��<:�@خ��I�� ���l`�n#+t!-���%�Ly��3�t�r�Mo�m]Pp�w'i ��]����po�8�o���e �f��D6��*U�94�e$�a���L�cN�����	
��#��0���(+�SC�Yy�{ޑ��r�K9�[�"a[�[��Kwz9~��c�}�N���pu�I4�Q��H� ����aM&��h�����L8S쌟�4-�q��-�R��U��!�I��aF�=�(c6���"i��h�f\�M.���R�ܑ�1��a��K��>B�I)�z�������x�}+�	�>����fېjM��L�;�T�N* J�7T&��*���Ё 6(kS�*�C�}�1m�QN�<�@�	c'��zzC�&c�}�s	�b�@�X�	���^�I6/�5.[�V)L��]�O%��<���n7._�5��:F}��H�ԑ�z�[�jE��O�C������
Y�^PoRy���WEʆ���x�� �D��$ʙFHE���uƮ[P�f�8��e8���7D����W��:S�iÒV�#���v��SM�j����v-��؃\�PyR�`�G�$K������C�!l����(A�M��_6��n�գ�K��!�,@ؗ�y_��-�^ԋ����*�(�I�{���9�p�9H����O�P���?0׳��W"�s���{�,�⊴g�l��;���������q�y�����^�ܪ1�,�F\�>�@������_kM9F��
�2�6\e#%�a"g�kb�Ŀ]t`��e.�1rNp�d��Bn�Z���\�u|=��,J�0�j���0�ۚ�>�QQ�����̱�����y�NNi/�Ԯ��P��/�;���Q�w^�����1�6 ���Fǔ����;�ā�U;0xb�T��u��0�U7�K��5Me�+Of"���Qun�6Q=�br�٭����v����c�^���ֱ>B(KkfZ&5�ԁ��Ij���3��m�3��"�
Pv�m*u@t�����t��K>GA��)�M�͚��Ҟs��H���cZ�GqP�
��o��c�>g@��/+ĴB��2Wc1V1'��t�H����s%��#�:�����?�n�nJ�~m�t�E�U�͚�AUQG�3ar�U�����S��y�4����-妑�0��p�({���ͳu(IU��z�:��2&�X>��f���1����ݠ��4[��f��՟P��4�0L�WK�LJ�Bӹ�]Ǝ�x���Q{�N�^PK�N��r���A�բ���U'8n�*��C��Dm�����u��:�����<��Nv�@��̨�������a�%a��v9����[�o�E�D���� �h��oF	�-������%�ua���\;�͙;��J���/x�#O�h�������zݯ@�i�g�e���� ���|I��*_^���"��2�ش/��P*�9�úHk����K��27/��q$$���� -����x.�b%�_���}��l��I	ά�$���X%�Q�)��EU�^E��f`�T�%�ب�WVI�,֊��/Y���?l����s��	����9�Ӛy;g���{p�m��s����f��i�$���wE=���s������T�a�B5PM���\��>c ���%R�l�G6�S[�c'
�=s�w�J"�9�m�G\��z����mߝ~37��-�;�����$Z#_]$qc�'�ag�=ݽ��۠�g �&�y�$3��%�\����úJz���(Tp.��"5��Ǝ[X��6�������1��2j�� �����wS��o��G5(?b?��['�i�H�.���*�BCB}�eX�x�j����쇱�nP�z�t$�FX��Q�3���Q ��B[���F�Gh��qߊ��%�����$���3:���}�S.��%��h�I���,�}\£m���L�W���R��&���%����PB"�A V�5��o#�d�s~�h�Br����q(�M�ܒ��IZ�lb&�Zv`��=
�l�`�8����~��[A��˴�����F�r�Q}�e��<�9b��x�E�ËU8/�e�\5�\�c�m:��Eҭsfh�Sӎ��PT����>�	�K������=��z�(I��Y�W�")���v��H/�u:�	1-�8��zU�Ew|���$��+�W���a�(��[=&��:]�	�p@���V��l��37)@� �bBS#������v�T��M}W�|G�K�_�����7T�GMo�gBL�{*u�э �x����P����Y�Yi�r�L}I�2�UE&�H����hw�2�"�hc4��(���;Bٸ>�����x��sl����1u����'�j���v�	�4LT��m����ڷA�������L�%5tpC'��������� �q����.7��0�(�|��c�4�X��˨1
��c�laÏ]�ݵV���~��#�x.�Z�fT��W?�X�Q@�BfdCӫ'Y�4ة���MQ��(
�VOJˇA����4�;�MP��[S�F>���%S3Nv��y���>�
5�Q:q!�Aa:���(	b>g� ��G����/�=u��C������N��U�����1!˒'��'Dv2����������e�į�W���!�F�o<�}�����u���ه��P^�|�鮌t%6���^��v�Kluo(rnV�L],���B@��OZ���R�ڂ���Eci���c+������Y0�T2�,@�jЖ@��NWm�������ׂU����PL�$i��^S�w[��I2��,�<���A~�(���MY�VFm"�����
�,Ӧd�I8�*Q��4�E|���������6�F^��o��_y�tA�}��dq�8<���Q��T�����[�(I�l���b��9����b���Vch���!�b�`�[VY�ߜT�
����E��i����xp�/0U%�e�C�K&-`C-i(d�R�cPa-^���p�E.�a!��ֻ�O֩.t9�e��;�D-�{u�P� 5zy��q�5Ӌ��Yr�g��uB��>�%��Rn�q��5u&����C�?�h���e#��?��{@�8�nu��HGB��&]�bT����y��$ڹ,u��N�l^���� �E&���%�D��- @G]uO@����x��sv�G���slc��]����\�g-A�~���6@Q�vp�j_����Y[/ڍ;� �И�i[�U�|7��]9}� �,G�s���!Y�Hv�e�J~��m��e������?� d���+�7B1�3�!4��B7�����ƦE�)���_���T��.��EQ̋5��B���u1^�>Xc³�骚�	���Ӎ� �,�΀�+�S��@?��	HkZ/|XvV4s�Ⱦ�e_�~m�C�z�N����A�8��#��$��/�S�X����8����zՉ�,1ܼFC��a"M��UK&�`D�l���2�4�+���F����7ڀ_��M��Y٩UZ�xyF�g_7s�s��Hh�A�C,[cƆqڳ[�>q�;�xX��S��W�Y���-����TY9��S�|�+��T$���4Ԟ��x����7߁���y�����D���u�q�J�N���ՕѼ����,��y����1}�G�,]�$E��k:���b-�	}��o[o�XR�=D��w��׾F����e�I8R��S%���Ή8y6�U` �Kۺ�P�o���+x��z��(� lK�1�x;�w�^q����㸴J+��7�Y�K�i_X$d�E�� CHiXH�c�.��8�M���WD\0�a�i��U���0k����M�ӅQVp��d�����[)�ĺW��Oy�eX��'��c�Ai�+^	���v�k�u={��0MH�����rέ1�A�U�(���7D9SK�$�q �p�ᙞ���?s�%1�IM-�`�덧)��=ѡ�*(���4M��5RP��ٽr������0�H+/B}h����$,#��8q�x,Qĉ�����n %���ӝX��ښӸ��M�1�g���$��m�p^_������T� �Lo��`~�J�g�wF���o����%~m��B� ~��j��.�f�u�0�d���	�PG��I��V�N���R��[E��{"�<'Z)'�~��֑|���6��2��\���y�7"�Ͼ�>�^4���X���,�ބ�l�7�+���8��`�~�]���=bG�0>�L�a��#ˑ��ܪ�����Ԁ��ڜ;[f"���Wy�J�
hDI�E�;Ym����ɉ�'0V��.�_Ȋ��B�'��J�����I��n SȳZ�K�bq�s��Y�T���l{y�ϝ
����4&������s�?v��U��ҚD���N8�� �,@xo�mPO$�ه�dh�4c���w�;�EU��1��53��%�Ŝ���K#Rt���4���̠t� !��e�Wq��Ge�y�@���\�o$�5Р@M]ٸ�ܹ�ɵf�� hC��P��ka�~p��L[����8�II��#���p:�zI��xo1�#���%Y��M-�p�A>�=f���ZR�,��X)�v�WǮ���>;���_�Wѣ�se����?HV�oQ��"�Zm�,���_�_�,�Łt��JrzY��O-�D��v6��y#�ri��U&���I�/U�ď�d���5�~��j��+�d�3�u0@л�����J�P�P�(,gv�6E����$�6
�>��KD�ehz��jYW/av��s;�E�+�_�� }<�Xj�V��lQn�?��DysZ�n�ɍ�S?��J�m�R%�w�)�4I������B!��{N�A
X$�	Z��gƅ�S�z��&�]�`�7���׺��fUԻ��Ž�o��5&��1��5��V@�Js���S!�*�j����C�b�s���Nÿ�0��r����R��T�F�]��i�8͆F��� ��/^]uB��Y��I؝;Z�[�%�?�3��ƕu�{�u�?�l�pNK�x�)ilϔ��<#�(�V@=e�`�!p�`�eF�����뗠m��q�re���Xrd�)T�xf��ի�ME&�ЖmCV]ÎC1}��fk�S�F<����Y�3 P1�\����]�����\[0�1�.�/깈mZ��ZS��#S�F�ӷ���m!@���q$m�%��'�����"�ѧ�	�c
N�"K��{���+�K����u�����R���c0��?���_���C�m��A�~�nS\� ��%b�!�p��#�0�VqQ��%�n}�_z��I�5�f{���5�_Я�i����n��>7]�ȵG�W��J���R;������A�-PVE�����Ӵ��տ�׏�V�׭�h����Gۚ>��'�cA~�u�⾘��m�ؙwM�~6և�.���oe���KC��O}�/�gH�/�� k�5�ɜ~�tޭg?��6�������Zs��-�b� �vM���3�~���OpqE���0�M,�l~�ѐ̬�C�@m(��8��RˑkԃSH�T/����`�!>����AӦ��W�m���~�&�\u^�U<�_x:���]�x�c��/�Iu�ױ
]m=,����m3/fƳ!b?����u���*]6�y~���l"���-����pawΌ���ъJOu�  u�90�����#>W�|��ߎ�θq�&YR�X�d\�&ᰓ�6�kn�i�����*
��F�9�Fv��tl M��mP�^�H��1[}�V�&���LN�C����7��@���&F��g����,�h�������@(����d2k���$�(���z��0�&�i�L�5�q��IuNzeu�)v�q� �G����#�G�4j�X$�nV��%n�!&A��!�q"��8ӆ�+�$����_���N_�
nO����)�&8�% ��yp��R6eQ�6�F���d�|$	�N*�Tڝ%Ԛ��<�R��~2��<빱�vx���(�M	=<X��-_�&3�y���q�x��� �����=�P7�D������t��2�|N�<���FR2�h����Z :S{�F��z�\"��'8!W�h|���R��8P�*z�#9'-ߗ�3w
��9/f��RZryG���Σ��6+4�[D$�,��$
�ϳj�ď���1��7 ��o��w�`�(X�/\��';��@�W�ǜ�k��|��+M�c�\������LuA����V����ٟ��آ�����tDA���D�GT�_0�X[�L#>�[ΨHp�w���e����"ޙ$�#B@�0����g+��^[1O�e���p�E��8ra���oA�1�eA�/"��_6o�DQ �op[����R�����l��fHS�5x\�]�$ +��z���;���g�&=]��+�I�VA�a����6r��Qf�d�Y��">Ut55\|~q�+8%�+;�u)���$K���+�u2ۄ��ɏ@��*���3�ynX�o&G�7R�r�?�߷~b<B���H��º)�}m�`�261<�9�$�8)!���w��0�ؓ�Dv�U��©(i)}�&����E��Ux�YH%I�A�ǥ˂��cs{����	߹S�m"��[|�J����låzR��$����sD�|4����s1�|��mu� �|OOjX�T:�j2�R�@!�&S�G�Ƶ�oÄ�3�w������)�O/�v�\����TXGGR�	4�e������Z��Bg�`��R��{d߲��ߦ�.��1�s���ƗR��[���S2�ҫ�^�_��t�p�`|8�J��t�f���b>��H��
�K'|G���ѽb��!�g�A��au;eeU�Q�+�y��pZX2_F�^]0����3�����s��F��T��3�i�9�ۀc�?��.Hp�A��\fv�iU%��.^{@.�UM��h3>QPw0��Y@D�dd1�5��O�[H���{�;D/Z���`�[w�b�-��5�)gX���x���a9��=����_�>�AO��Ϫ����G!|@��q����f'�i
y�A�n:bz1�T�,IA���;c�G[r4�ǥ3���9ȉ�n'��k�5-�$�f�����cʪ����wM^{yo����ۙ}ٝ>:��|v=P��\G'�MB�*��W+]�g8Z�̊�'���M���4$�A>�k�)#�1D�h�`6�8� /�If̿8 Ͷ^i�6��n;~1�2IlC�_D7�B+ѫM�M�9���n;=�υD ���#�(I!pbnkK:��(���-h�z�h=��T�$��L"�R.D���VJ�k�!v���z�[;� �]�$*��pOz����f�?�ڥ00�Z�Y�|sg�h�XD�x�����mX%�#R��)�X��@�����P�L������4�6�vn2��J���X��P�
kG$�W�:+���~6����$R�qX}C��8� ѦO��<����q�,�;��	|2L�Tb��y4
hU�z�����+r+:�:�[�|d��m��l%��ǵ���0�o:ԄV*��f^�ȶ
��9�Ў+�F��3b�?z���.�%�x���l/�V'`��q��������ܷds-��B����u}3��Y���.�������Z$8���r,@�F���qo��WD�������fk����&D��B~�5O�j]�;��:�*$�̕�!��x���B��`]gn��9�\���3"� �@��h���h�ZS�=�X�.h	��W�#��ET��R�n�
�X���q�J�'I��O
c;�9�3��}v5@������p��2�} T!���/��8~,[�è�P�pϷ�N0)�r6d:=ǧ�9Gj�)�$�2"�t{7��ؔn ��������GJ���T����d|~>�]�kq����:�3v�o9�W�e9��������@����U��pfƣ�E�9�Z�a��~d��Ŷg[�V�Ք�s����o�(I+Y��/.z��5t\����p{�mϑ�;I�'˓=k���k�tR�'�q&.$�i�Io�4�Y��:`^☌hJ_L�;�I��|�[�8tyE�Ȼzѱ��俟�MGl�Ȑ�a�}�&���ӰpPX���W���c�-oeq1�K`SOvVңc�B���'�=��s�l����_`%*E6Fh{�d��6�Y[gB4��^WL�؀��׉-��vx��jZ�a��(�������쯞���u�>ՠ�)���KA��⾆H���\2H�64S�a&�.(��!x F7H�^O�!�}��8��t��d��ٷ#-̗��s7
|�����q�u�R�S)Y���_����#���4�·E$f7��ݿ��^����I�z�r0ZoAj&� ܆5d�4*�u��s�f�Y�7_G3�/�6!9�Х�R[�8�韭3����⽻o�C��u2}}N�_��rӦ>�݉��[��v�g����w�A:�T�F��|-.s��'�LC��Z�B�&#U�3P�őM���|-~��πF�
�?��\:� ��*���������9��&��Qãj[*7}$�q����ڏȾ��{תe�P�� ϕW*0I����T	s��r��B+ 5Q��`����xV��B�C��ݨ���{m��"��<YD��jQ@u�����]*�%b�(�����a;��7
ŉ�b�:�%�5d�؈EMw�~�(��Gg�0�.B��M΍���l� H7����?��x�
ː�����s������ ��3YJO� �����`�8 y��8X]�y#pj@����z��#��P<�լ�j����� �ѳ�,����|�����kU׾M+MO�p@s�֢�b�t�	����k����*j�Y�5�����t�n�зH*M^s�<��ﰲ�+m���	��/����)\G���6S
g9g`��އ��R�� �#��7cg�myTD��a�Iq��:pM	�8p߻FY����6�P���1
eү'��5�M�)J6�&ZTt����S��x^���������*!C(s#�����zc;��I'®I`�-� ��x{��~r,����5���Z�����l�}4��S�P �}o��L:��4b��Q���.M��ZT��#���k�6��G� ����tw������4xʌI�6�,u�C��L(�*�	A���l3\���\J�aɟɺAB>���v�,����s�i�&�"��F���Ew�	��آ[C�S� ���w$��:�7��chϻq�f#r�ݐi'��R"�y��3��C �8EL� �h.��%�V�nح�7�$'�h_	í���䱧�(~��z[�[A4�ɱ��0���c��P���� �D+����U8*�C;�������,��f
�*�T(�@��6dR7�x^�TQ2kb-V4���B�l\�э����<��\��<��
�?�{��=t%��RC@����>�O
�����!���ߏQ��p`R򟞔>��74�{��4�c��-�l����uqE^�ᨪ���Ɉj<��"��^��O-+ҧ�'Vi@�:�/�)�t}���F����?�E'O�
.�������!Te�k_6�R�}	O��ccZ	�=�7`����­7
6]��XH��v+&S��Td�C����ᘶX�M��}�B�Y�Z��Y
e
Fw
�0ei��j�R�z��4�KT�T��v>k�O����s�]���2(�U����i3D4�$�8����}^����ݜ*�w�Ɋ�v�du,a~��V�$�'1)C��#�nT]��(F�԰���A�&D�C~�aZ�������u%�-fK�"�]%�SN�(Y��f�9U�-#l4ð��eݣ`��������I��� *��c�G�?7:�bP��	��)*���[��@�5W�b*��o^�R�zE��e�8�C
��w���v8�Ւ��se+�<n��?����^���:�	xnB-��L<���hs��UyZ$-yehp�JJr�����&"8��)7C*_�ns+��iy�k-Y�ɱA�����¹��YA&؟��� ��")R�t2~�g�pj�ShL����}Jy��m=�u�)d�T4� ��5R��v�*w�>L]p���}�ƌ���&�D�"�dB��5@Zb��MjB���M�#n��n�%97�uE!av�\s_ҿ[2Q��p�u)�l�z��q��#������j��٬ۇ�F}�+��%	<���A���1�l���^�^���l��j���ǆ;�ig�����Y�چ[��BY^+w��� ��0ѻ+�w�ŞG�� �f���[i���tiْ1af8�{l�2�5���P�b`�ɯ� \�*Z���a�/Hk��5������I�L�ʦSfs^b�t��;��S�J���KEO�'���'�D�M몝��n2�HN5��t��x�5Ƕ�𳬽t�o��rd�F���"�����A�V�ƥ��C#�Ð�6��~�K٧�v�	��BDD��C1�Z4�נ��Eў���P��+._�0[f5h�MѸ,2�}��e�&��Sc�"1���B�ڑ��=9�ᑦ!�e�mHqՓ�bm�f'�p�T�:�-���\����+��n�xl��������&��g?������I"o_�~ģ�P�Rb�e�}�����xƱC����<��Irf�g�-&��4�@~h��/-9���X^��i�b�����˫чxD;��4G̶(���ᮯXI8
Sb9�-��*�\� ��E,�{�R��[���
,����+��m�	ӆ^�)D88l�p������' ��e2�����KV���r'��%� ���ы�X*%�EE_["��[ّ�F�I3D(��|�C�Ћ��9�G,�  ������ [R��Y�����uE��!9���Ȏ�2%�0\��8�N�����B �ߵt����ANyZV��ֶ�!D&����eM�YN�����Ҙ������iK���*_��I��$1���o5�1v/M�3S�I��v}G�f��1�̨xee�������J&�����J=�{�Il���X��l��\Qhl���YkR|F�Y�iDt��b�}�f}g�(v��?�T�>��nCf'\�_8�giӈ��R;�5�fZ?j���ꭋQY�u&�� U�v�9����h����T�3b=f����Z%�aC�Xc���;���2��3��XĮ����R&��!k�\u��m
X��\�(�q����rB�T�!�&���+0��[^k�1�	��"n#(�3��&�z����;�Y�,h{�SVfrmv6������4/d�d'S��ޮˆ�6��Ν��n��4b���!�r��˛�5�J������b7����&����
�#-��5hg,�
hc�����:'W
Ҧ������r�շ��hC��h�0�#��qp�yU�yޤ��	VN�KN�i�&����2-�����͚�j��w�������E�ߩAܴ�1�R�j�e� '2�t*�F�C�̃u����ݛ�C2%`��Oqܔ����+K#d�~�'��AK�2W�����QY���P݄]
}_�-L�r��;��E��y0�i	�~������3��aXћ�i��A�)�ڛg��r1��d��0re�uP���1ж���u�7�8є,�+�5tx��>�?�����M�h��n-!H�����|/��� Tf�䪲2;���v�t�W��"5���Fi:�Q�)�82�r�4z9��z�S�U*��)A~^���'��Q��.�����7�H\�Ga��ɥ�:����aPs�|��v%3�N�=�W��-xz�P�_�]���#����V]g�0��?�a��Q|Z%l�`�1��B�A~s`2M�=���5X� �Y[MW���(�n�9�CJ��+��mcK�P�O�ۯ�0E��6����,҉�m���ǖ�ĺ`�j�"$I)e�j��g�ߓAjk!��Ȑ�?�Q���A���[���ڐs�����3�{�f@�ëC���{��u9��8�8�@<�~t����A8<�I���'�j�%��_�~�����i-n�x��@�{@|����+mD����X[V�Q,����r�1x�����h�WHT��g��'97�NVK�q���+<��#]��A�u�^�$���+��ۇ�ȣIu֟�����3����
�ߝ�	ڎ+�7����¿���v��6��O)���*a'~�U�}�[�3�7W�#�o�%�F��?��O^X�^�(���9"�#�Kєw�����YBW�=�r�Xt�v��̅��y��	����[	Jwb�*�l|����9�嶳���s��\҂��R(����{��p���Z��M��M�z�׌?�s��٢Q��m����u�B� +�3�ײ��=��o�Tdm�K��e�֢��
�H�Ȥ��0!E�'G�JD��k�7��R�ؠ�sm轩RP���?����J|�$ű:(���n�ǬnKF��C�c��m��C���%z��uQ���]�4�o6��x�W���� �� ��0h��:�<��(}ꊪf�ظ1�Z�� O��G�7�������D�o�0�)9�n Z�le�t+���?r����aH8f"���ϖ�9+���k{��"X��>6�j��*��2#��#�b�M��a�w=2�2��)^��d�vy#��Ig�{�0��O��ً?�η�>��r�;A�$6���z��p���	�v���d�YV�X�"k,^��G sWR"�&�w�>Vko\FdEx�mY�h��B��O���>�G+�՞����{��/�z�H�48���PQh4 {��@�����q��+���vr(bB���%/ţi9�b�=9^����\����%��j%F�"{����ǟ�5�>2�����{{���EP�7\6�����~��Z.rA��}�!�u)�NB�'~�2�z�{^��М.�1�tnN`��h���f�߻�B1�v��dQ�X�*]��z>�mR4��`����k�L~,w�;b�"��y2S���o��l��޸z�t�]ź��tQ�e�o֟�m��*�r���p�/�����+-pຨ��6Gδ��#��_l��
�4)�RK����;�_���p�!�w�0X�m�{A�M�����r�D���3%�o6%5=M������ ��L)��'WmQ�\K�7�pf?��!�33bu$�}�����Ϝ��@�ye ?i��ŝ�=bE<�jQ:��H ����u20��c�",���т������w���u��beg�е|B���s_���b
NB�\�?`O,�P��PI��ȭk� �C2Q��t������CCi#�
<�]��^<��Pi1��gk�k��.�<tEut;>+EVc��Pw;�R�b�Q�K��Z�������00�@a!�M!��8�@U�h�=�T�'k�~��}�v��7]�����Z�o�"�}qN�{��1Q�m:eϺV���*:����W�7�6�,��mvך�SA���b��V�ЃMV,v4��P�Zג�c�����m�<����Ҥ�����ȨMBE�@-���?��m��A�>+6%���Vg�bBiv����x@bo�h�W�����9`ɼ5�e��̝��Dk>X�Մ(�Ш}�j ��y	­8u=���M�c���9>�UΆ�����5$}sj��q%��XiWU��=�q�#�:����[�yw��)#��R�:W���*g��8��P[l}���u��G����f��$4�pj��2Ph0�琿7���]�4�N(�38�r�f��j���� Ou��;�{
D>*5?��d=�*?]�`A��T�vIe�6�=%
STٜ!�7��70��U��CDE�t�)(.�f��c�W"�l��m�c/���;�]Z��Q��*�u��%֪�.f����T쀤bc�Loc͹��p�p��P	�RfaJƞC��T�#��/{�T	h��f�y�7����r{q?x���"w��s'ʎ���A|�zk�}�a��D��^�=����<�p� �{	`��R8�T��s{�(�Z	l�qe}�i �0����(�hG����*�괘M�/�$�2WP!1���~�<�m�G%̗�?3�zd���Q��U�m;���m_����n���*:�kw��q��1ʡZ�Q��� u���+����<&��h��f�ήiF�|��������D�+�Fu�e��UV:6��A�>4�p����'U�в(3�_�"����/� 9wDT�5E�z?�$�hb�k_���CzZ}a�� �c�<����P�N-s��E�$��Z���zEd�T�e(ƒ��.��x%X��_��%j;!tgq'�ȇ��.4���,!5����y,4�Սo&�_��P���*̴�-^��b�J��i���$?��!�!<!���M�>��9�f��\鲿��݁�-�?h��y�P������q%}������0mC����w��gV%��m��<$�g�`�yœ�`2%����Fh�e�h_�@�宾��W�~B��~ڄ���=$}-	�v*���4�X��4�_׵��`�PB]�hф7�<���U�Ij��%t_Vk|=��%1�m���TW���L`� ���' ��:^��l!�9
u�����L�B��Ü!-	%�мЉ^�@�IrB�1�����Z�4���W<U�MT���ӝ���-`�=�a�W6t�K!p� ��SV�~�E�l�r\Q4�́Q��:.�9�Nڈ
PE2:��h�g�pS}�46���Ư�Dm3��=�$-r���N��ղ���)W#S1P���6��[���I���rNb�rK�e��6ߞ�b���z{��`����ؙV�κ�|1���w>�4w�sh��T�	�1�3!>���o�/ۀ�Pӈ`�-:we"�ɏ���6����GB��m5R=c��i,ե��媁�hL�kvw0B�o�X�6�q��D��|�;g�b���V|��C�v&z�՝�ml�cY�i��l{��)C����n��o�Ū�QX�����9���g����׏E����;��d��'��.��چL�u||�(��ʺwv �c��ޘ�wv^c������;�B�e�P�;��`�]򜷛��;���ΩXнo/j�)���/�k0��)�z�i.�8�J�ہ�U�*I- F�=�B�K/'�i��B@ڽ{���+�ě7�7c^�>���]���4��� �T0���Q>B������-�˿�6�tJ�a�[�>�#���P�g�x$6ϖo��e.o#�N����o�
g�,���m���B�B�i�l�t�ߎ͓���uxH2IS�����0�yG	{�մ��6a��,��G�e��'L\hf����nV�d�9'�>����^Fg~�5��+#sf�HD�������05���BA��9c�q�K�w�8�u���d ���v	� ^����\|�o�Ȋ&�~���X�0�#�ykt:
	o�n#��sG��$tZ�سx� ��Tc#��0 ���}���2�T����7�(0����$��#��������c��u�)�Fdٜ`0<�DQB�7k�	j�Z����F[D��X�$�W0���t�#�/}���K����ʃa����-�!.�ΐ��@�6x��8R%Um�Ly�2{������y��b�C�7����Q+���٩�x��1w���a:���k�_��R@Ƹ��x=��<$VҼ��l���z�;��\E�F�ϭ=�׾�e��D�R����G�Qz�W���ѥZ�i��v��-Ɋm1]G}�lE��/oN�-�6/;��{�ۮ��kw�
��ҷ�J�������[XN�{�t3�d|O�~T�m8���'ѶV?��q��b���b���=d�`ˮ ���o�e�.T�hX!��l6���
���d;i��T�<mm!�U�K���Ӽ �@�/�� �<*_$��ԅ�,�K?�����Z*4擸��Q������bd����,�+Np�q��W���+ֵ�3�1��!��.E��A��[S���4no����lj��|,qZ���vM�-.�{�PuW;�6�s�s��f��q(�QGz��Rf�]�?�D�9ߨ]�B��L�E?ξ�$��n�8����|�xm,el7/�1[��޻l/4!8���]��֪U-"���2�J�ׯ��L'�m�?�ZV|%���(��W��M_�%v�7bT����7�0�Ah1�ME�}'�F�����H��K���C�f)������)/���{��r�0���k2[��np���$=��53���	�eQ*����TM;p>ȚPM`�����-]�Jt���:[(�O������L<zO-!էt.�JBz\-ģN�8g:���^W��"��`����`�}�?-�p)#���6����M�M>�#������@
��'&�z����c]Wn�y8�7:�J��q��v<XC���τ�BF�Cm}k���C�a1����x_9��O6��]��=���
�����"�F�M�����YA|twZ ~�t�>���U��	v�X&)ȡ�����S��Cǭy��pȿ�L^�v�RT5f9��4�0	���kĒ�z�k��;۴�����
��Y���G"o^����C�M͗W����K��א�P�l(�7��[Q�kp��k�Qla�WA�����U�!����Ns�;�)δ>a=߯�_�f)�y��N�3�Ъx�g�p�
�;��uy�(��D�K4�8�xT5�k��top�f�r.������A
ւ�«�������G
��^����o�\/����^�pǼ�+>�D�d����X���G'=:��5��@��pC����mSf�ړ+;�����|�uH�=n���u沗 �E��[18����J0�b�<��To�X��M�$c����lp�#�^B�j�����Yn�jc�x�42U�LP9QS����}	a����/Ċ��3g@��-��dCt��|}A,]^I�a�G��&Q1֞��������ڗ`7�3V���7��J��:�K�8�ז�:��~��6�ь"��y鵸�VIY<2.���9� �E�d{���.�Y��$�zJ@=~ع���� ����^�;�p��r�ы���S�)��Y�e�:.E���̩Xz�1f%CCPj�lG��Sq��h��� �1�$��k��ގ��@��p���ų<��[dYN��7�y���+��u�(�o(&]�^^�A$834��5����tAZ*��Ou�85��%����.����p��[�i ��>g�Z�L/�.DU��n�|�]σ�=��[��G�rLPq#ʚh% z��U�0d��Z2�j�`�P����*�$S[2��D�yF�<ȕv����h�������'ۂ�s�V4�e^T[HI''�e�jtt�aу��|Ą�y+j�S[��&b������YƑ�u(;���X0��l/-!��za�/�xx7�$�����E�;����3���<���[�e4?�ǿi�H?{�hTP�wO3�r�Ә�;�58\���0�d���9F�~r�~�͉�zcK�2���Z�:���x��|e:��4w�)��'�~k�2��o�S���9M5�Ȫҏ���x�B{�qҗ� ΖΧ�A?��nW����pD��?�"��X���i!� �My��&�:$��A�Ρ�u+0�1^Y �z���� o$WX1��g',�<�����S3��u䪦���BD�q�C�=��M&o1��j����nJ�@����X����u?�+�i�Pܡq0oE�d1I�����-!`d�;CnC�g����j'�dm�.{�'��j�����I6���c��(����	��>��P�xP�?5����;����Wfp>o�����:2V�h���OI(���wX�+��+� ��E(�;�$���G6��N�	�}I��pI����@��e���'-#E�P�ʂ�b�{�ɹ���$����M`�	��8�{�,�L_�U��H��~Ɯ�x�5ׂJ���_x.�ϕ	5�s�gݽ��*:�9mDE��s^��&L�E9���&e6��s��#�!��n#�J�m޿�	�����=�_ѵ�4 G���\{a@	�}NG8�#E��.!(	���V)`�$�*>V�:Aȇ6e��(h$ኄd�4#��/���!��\�t��V7<N�����2��xMG�9� RA�o�B*���op��s�H3�a�V+�o%�t~
�Ӑ�׃7����Y��v:��Cr�9�BkQB�m3�LY#�=�J�e�e��R5�ڧ�W��0����6�T��`9�-뉊f_��@}��������)�&q_j��0�$oO���b���E�g9+�O��,�)i@��kg��PY"ʙ4���i�+�%�~2�}��Ў�ZK���$�7t�I ��&���rp+e#l��T}���:��Z����s��4�S���C�(��~�EO���R�]\�|x:��t�َ�!8�_oM|�G㮙Je3��k���Z� 1~:r]��M'�Yj��X5�4�� �CTK%'v�gw�Vy��Q�^�!b	��*ɂ;� �c.d2r׈��w�6.$;�lwȁ�䷄�1X�iͽE{��A=�����[�Zo�S\(z�îQdR5�6�1D�����td�j5��8��F�F��am4��{��632��2AaGt�Z�.���A<u�����]��68�m/��7��t� ��\�èt�9�Tq*ϝr��F��+�vm^����)����@�r|c��9�7W�����^"D�׭3���)C����bs\G!7,����,'_���s��Si��l|���}C�[��Ȓ4��Ԍ��c�O;��M=N���p��ߖgj�W<t�pG��\܁��j�@��NdO���DX\6���W���5$� �A;͡o��L(4FD�